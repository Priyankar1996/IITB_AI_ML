-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity sendOutput is -- 
  generic (tag_length : integer); 
  port ( -- 
    size : in  std_logic_vector(31 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
    zeropad_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity sendOutput;
architecture sendOutput_arch of sendOutput is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal size_buffer :  std_logic_vector(31 downto 0);
  signal size_update_enable: Boolean;
  -- output port buffer signals
  signal sendOutput_CP_26_start: Boolean;
  signal sendOutput_CP_26_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal if_stmt_42_branch_req_0 : boolean;
  signal if_stmt_42_branch_ack_1 : boolean;
  signal if_stmt_42_branch_ack_0 : boolean;
  signal type_cast_51_inst_req_0 : boolean;
  signal type_cast_51_inst_ack_0 : boolean;
  signal type_cast_51_inst_req_1 : boolean;
  signal type_cast_51_inst_ack_1 : boolean;
  signal array_obj_ref_67_index_offset_req_0 : boolean;
  signal array_obj_ref_67_index_offset_ack_0 : boolean;
  signal array_obj_ref_67_index_offset_req_1 : boolean;
  signal array_obj_ref_67_index_offset_ack_1 : boolean;
  signal addr_of_68_final_reg_req_0 : boolean;
  signal addr_of_68_final_reg_ack_0 : boolean;
  signal addr_of_68_final_reg_req_1 : boolean;
  signal addr_of_68_final_reg_ack_1 : boolean;
  signal ptr_deref_72_load_0_req_0 : boolean;
  signal ptr_deref_72_load_0_ack_0 : boolean;
  signal ptr_deref_72_load_0_req_1 : boolean;
  signal ptr_deref_72_load_0_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_166_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_166_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_166_inst_req_1 : boolean;
  signal type_cast_76_inst_req_0 : boolean;
  signal type_cast_76_inst_ack_0 : boolean;
  signal type_cast_76_inst_req_1 : boolean;
  signal type_cast_76_inst_ack_1 : boolean;
  signal type_cast_86_inst_req_0 : boolean;
  signal type_cast_86_inst_ack_0 : boolean;
  signal type_cast_86_inst_req_1 : boolean;
  signal type_cast_86_inst_ack_1 : boolean;
  signal type_cast_96_inst_req_0 : boolean;
  signal type_cast_96_inst_ack_0 : boolean;
  signal type_cast_96_inst_req_1 : boolean;
  signal type_cast_96_inst_ack_1 : boolean;
  signal type_cast_106_inst_req_0 : boolean;
  signal type_cast_106_inst_ack_0 : boolean;
  signal type_cast_106_inst_req_1 : boolean;
  signal type_cast_106_inst_ack_1 : boolean;
  signal type_cast_116_inst_req_0 : boolean;
  signal type_cast_116_inst_ack_0 : boolean;
  signal type_cast_116_inst_req_1 : boolean;
  signal type_cast_116_inst_ack_1 : boolean;
  signal type_cast_126_inst_req_0 : boolean;
  signal type_cast_126_inst_ack_0 : boolean;
  signal type_cast_126_inst_req_1 : boolean;
  signal type_cast_126_inst_ack_1 : boolean;
  signal type_cast_136_inst_req_0 : boolean;
  signal type_cast_136_inst_ack_0 : boolean;
  signal type_cast_136_inst_req_1 : boolean;
  signal type_cast_136_inst_ack_1 : boolean;
  signal type_cast_146_inst_req_0 : boolean;
  signal type_cast_146_inst_ack_0 : boolean;
  signal type_cast_146_inst_req_1 : boolean;
  signal type_cast_146_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_148_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_148_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_148_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_148_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_151_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_151_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_151_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_151_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_154_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_154_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_154_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_154_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_157_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_157_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_157_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_157_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_160_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_160_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_160_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_160_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_163_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_163_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_163_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_163_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_166_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_169_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_169_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_169_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_169_inst_ack_1 : boolean;
  signal if_stmt_183_branch_req_0 : boolean;
  signal if_stmt_183_branch_ack_1 : boolean;
  signal if_stmt_183_branch_ack_0 : boolean;
  signal phi_stmt_55_req_1 : boolean;
  signal type_cast_58_inst_req_0 : boolean;
  signal type_cast_58_inst_ack_0 : boolean;
  signal type_cast_58_inst_req_1 : boolean;
  signal type_cast_58_inst_ack_1 : boolean;
  signal phi_stmt_55_req_0 : boolean;
  signal phi_stmt_55_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "sendOutput_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 32) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= size;
  size_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(tag_length + 31 downto 32) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 31 downto 32);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  sendOutput_CP_26_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "sendOutput_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendOutput_CP_26_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sendOutput_CP_26_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendOutput_CP_26_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  sendOutput_CP_26: Block -- control-path 
    signal sendOutput_CP_26_elements: BooleanArray(59 downto 0);
    -- 
  begin -- 
    sendOutput_CP_26_elements(0) <= sendOutput_CP_26_start;
    sendOutput_CP_26_symbol <= sendOutput_CP_26_elements(59);
    -- CP-element group 0:  branch  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (15) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_22/$entry
      -- CP-element group 0: 	 branch_block_stmt_22/branch_block_stmt_22__entry__
      -- CP-element group 0: 	 branch_block_stmt_22/assign_stmt_32_to_assign_stmt_41__entry__
      -- CP-element group 0: 	 branch_block_stmt_22/assign_stmt_32_to_assign_stmt_41__exit__
      -- CP-element group 0: 	 branch_block_stmt_22/if_stmt_42__entry__
      -- CP-element group 0: 	 branch_block_stmt_22/assign_stmt_32_to_assign_stmt_41/$entry
      -- CP-element group 0: 	 branch_block_stmt_22/assign_stmt_32_to_assign_stmt_41/$exit
      -- CP-element group 0: 	 branch_block_stmt_22/if_stmt_42_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_22/if_stmt_42_eval_test/$entry
      -- CP-element group 0: 	 branch_block_stmt_22/if_stmt_42_eval_test/$exit
      -- CP-element group 0: 	 branch_block_stmt_22/if_stmt_42_eval_test/branch_req
      -- CP-element group 0: 	 branch_block_stmt_22/R_cmp68_43_place
      -- CP-element group 0: 	 branch_block_stmt_22/if_stmt_42_if_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_22/if_stmt_42_else_link/$entry
      -- 
    branch_req_64_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_64_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => if_stmt_42_branch_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	4 
    -- CP-element group 1: 	3 
    -- CP-element group 1:  members (18) 
      -- CP-element group 1: 	 branch_block_stmt_22/assign_stmt_52/$entry
      -- CP-element group 1: 	 branch_block_stmt_22/assign_stmt_52/type_cast_51_sample_start_
      -- CP-element group 1: 	 branch_block_stmt_22/merge_stmt_48__exit__
      -- CP-element group 1: 	 branch_block_stmt_22/assign_stmt_52__entry__
      -- CP-element group 1: 	 branch_block_stmt_22/if_stmt_42_if_link/$exit
      -- CP-element group 1: 	 branch_block_stmt_22/if_stmt_42_if_link/if_choice_transition
      -- CP-element group 1: 	 branch_block_stmt_22/entry_bbx_xnph
      -- CP-element group 1: 	 branch_block_stmt_22/assign_stmt_52/type_cast_51_update_start_
      -- CP-element group 1: 	 branch_block_stmt_22/assign_stmt_52/type_cast_51_Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_22/assign_stmt_52/type_cast_51_Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_22/assign_stmt_52/type_cast_51_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_22/assign_stmt_52/type_cast_51_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_22/entry_bbx_xnph_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_22/entry_bbx_xnph_PhiReq/$exit
      -- CP-element group 1: 	 branch_block_stmt_22/merge_stmt_48_PhiReqMerge
      -- CP-element group 1: 	 branch_block_stmt_22/merge_stmt_48_PhiAck/$entry
      -- CP-element group 1: 	 branch_block_stmt_22/merge_stmt_48_PhiAck/$exit
      -- CP-element group 1: 	 branch_block_stmt_22/merge_stmt_48_PhiAck/dummy
      -- 
    if_choice_transition_69_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_42_branch_ack_1, ack => sendOutput_CP_26_elements(1)); -- 
    rr_86_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_86_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(1), ack => type_cast_51_inst_req_0); -- 
    cr_91_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_91_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(1), ack => type_cast_51_inst_req_1); -- 
    -- CP-element group 2:  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	59 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 branch_block_stmt_22/if_stmt_42_else_link/$exit
      -- CP-element group 2: 	 branch_block_stmt_22/if_stmt_42_else_link/else_choice_transition
      -- CP-element group 2: 	 branch_block_stmt_22/entry_forx_xend
      -- CP-element group 2: 	 branch_block_stmt_22/entry_forx_xend_PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_22/entry_forx_xend_PhiReq/$exit
      -- 
    else_choice_transition_73_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_42_branch_ack_0, ack => sendOutput_CP_26_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	1 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_22/assign_stmt_52/type_cast_51_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_22/assign_stmt_52/type_cast_51_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_22/assign_stmt_52/type_cast_51_Sample/ra
      -- 
    ra_87_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_51_inst_ack_0, ack => sendOutput_CP_26_elements(3)); -- 
    -- CP-element group 4:  transition  place  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	1 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	53 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_22/assign_stmt_52/$exit
      -- CP-element group 4: 	 branch_block_stmt_22/assign_stmt_52__exit__
      -- CP-element group 4: 	 branch_block_stmt_22/bbx_xnph_forx_xbody
      -- CP-element group 4: 	 branch_block_stmt_22/assign_stmt_52/type_cast_51_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_22/assign_stmt_52/type_cast_51_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_22/assign_stmt_52/type_cast_51_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_22/bbx_xnph_forx_xbody_PhiReq/$entry
      -- CP-element group 4: 	 branch_block_stmt_22/bbx_xnph_forx_xbody_PhiReq/phi_stmt_55/$entry
      -- CP-element group 4: 	 branch_block_stmt_22/bbx_xnph_forx_xbody_PhiReq/phi_stmt_55/phi_stmt_55_sources/$entry
      -- 
    ca_92_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_51_inst_ack_1, ack => sendOutput_CP_26_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	58 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	50 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/array_obj_ref_67_final_index_sum_regn_sample_complete
      -- CP-element group 5: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/array_obj_ref_67_final_index_sum_regn_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/array_obj_ref_67_final_index_sum_regn_Sample/ack
      -- 
    ack_121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_67_index_offset_ack_0, ack => sendOutput_CP_26_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	58 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (11) 
      -- CP-element group 6: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/addr_of_68_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/array_obj_ref_67_root_address_calculated
      -- CP-element group 6: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/array_obj_ref_67_offset_calculated
      -- CP-element group 6: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/array_obj_ref_67_final_index_sum_regn_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/array_obj_ref_67_final_index_sum_regn_Update/ack
      -- CP-element group 6: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/array_obj_ref_67_base_plus_offset/$entry
      -- CP-element group 6: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/array_obj_ref_67_base_plus_offset/$exit
      -- CP-element group 6: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/array_obj_ref_67_base_plus_offset/sum_rename_req
      -- CP-element group 6: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/array_obj_ref_67_base_plus_offset/sum_rename_ack
      -- CP-element group 6: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/addr_of_68_request/$entry
      -- CP-element group 6: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/addr_of_68_request/req
      -- 
    ack_126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_67_index_offset_ack_1, ack => sendOutput_CP_26_elements(6)); -- 
    req_135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(6), ack => addr_of_68_final_reg_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/addr_of_68_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/addr_of_68_request/$exit
      -- CP-element group 7: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/addr_of_68_request/ack
      -- 
    ack_136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_68_final_reg_ack_0, ack => sendOutput_CP_26_elements(7)); -- 
    -- CP-element group 8:  join  fork  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	58 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (24) 
      -- CP-element group 8: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/addr_of_68_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/addr_of_68_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/addr_of_68_complete/ack
      -- CP-element group 8: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/ptr_deref_72_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/ptr_deref_72_base_address_calculated
      -- CP-element group 8: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/ptr_deref_72_word_address_calculated
      -- CP-element group 8: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/ptr_deref_72_root_address_calculated
      -- CP-element group 8: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/ptr_deref_72_base_address_resized
      -- CP-element group 8: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/ptr_deref_72_base_addr_resize/$entry
      -- CP-element group 8: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/ptr_deref_72_base_addr_resize/$exit
      -- CP-element group 8: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/ptr_deref_72_base_addr_resize/base_resize_req
      -- CP-element group 8: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/ptr_deref_72_base_addr_resize/base_resize_ack
      -- CP-element group 8: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/ptr_deref_72_base_plus_offset/$entry
      -- CP-element group 8: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/ptr_deref_72_base_plus_offset/$exit
      -- CP-element group 8: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/ptr_deref_72_base_plus_offset/sum_rename_req
      -- CP-element group 8: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/ptr_deref_72_base_plus_offset/sum_rename_ack
      -- CP-element group 8: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/ptr_deref_72_word_addrgen/$entry
      -- CP-element group 8: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/ptr_deref_72_word_addrgen/$exit
      -- CP-element group 8: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/ptr_deref_72_word_addrgen/root_register_req
      -- CP-element group 8: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/ptr_deref_72_word_addrgen/root_register_ack
      -- CP-element group 8: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/ptr_deref_72_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/ptr_deref_72_Sample/word_access_start/$entry
      -- CP-element group 8: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/ptr_deref_72_Sample/word_access_start/word_0/$entry
      -- CP-element group 8: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/ptr_deref_72_Sample/word_access_start/word_0/rr
      -- 
    ack_141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_68_final_reg_ack_1, ack => sendOutput_CP_26_elements(8)); -- 
    rr_174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(8), ack => ptr_deref_72_load_0_req_0); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/ptr_deref_72_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/ptr_deref_72_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/ptr_deref_72_Sample/word_access_start/$exit
      -- CP-element group 9: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/ptr_deref_72_Sample/word_access_start/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/ptr_deref_72_Sample/word_access_start/word_0/ra
      -- 
    ra_175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_72_load_0_ack_0, ack => sendOutput_CP_26_elements(9)); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	58 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	23 
    -- CP-element group 10: 	17 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	19 
    -- CP-element group 10: 	21 
    -- CP-element group 10: 	15 
    -- CP-element group 10: 	13 
    -- CP-element group 10: 	25 
    -- CP-element group 10:  members (33) 
      -- CP-element group 10: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_76_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/ptr_deref_72_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/ptr_deref_72_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/ptr_deref_72_Update/word_access_complete/$exit
      -- CP-element group 10: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/ptr_deref_72_Update/word_access_complete/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/ptr_deref_72_Update/word_access_complete/word_0/ca
      -- CP-element group 10: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/ptr_deref_72_Update/ptr_deref_72_Merge/$entry
      -- CP-element group 10: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/ptr_deref_72_Update/ptr_deref_72_Merge/$exit
      -- CP-element group 10: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/ptr_deref_72_Update/ptr_deref_72_Merge/merge_req
      -- CP-element group 10: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/ptr_deref_72_Update/ptr_deref_72_Merge/merge_ack
      -- CP-element group 10: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_76_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_76_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_86_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_86_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_86_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_96_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_96_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_96_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_106_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_106_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_106_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_116_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_116_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_116_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_126_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_126_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_126_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_136_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_136_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_136_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_146_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_146_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_146_Sample/rr
      -- 
    ca_186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_72_load_0_ack_1, ack => sendOutput_CP_26_elements(10)); -- 
    rr_213_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_213_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(10), ack => type_cast_86_inst_req_0); -- 
    rr_283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(10), ack => type_cast_136_inst_req_0); -- 
    rr_241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(10), ack => type_cast_106_inst_req_0); -- 
    rr_255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(10), ack => type_cast_116_inst_req_0); -- 
    rr_199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(10), ack => type_cast_76_inst_req_0); -- 
    rr_269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(10), ack => type_cast_126_inst_req_0); -- 
    rr_297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(10), ack => type_cast_146_inst_req_0); -- 
    rr_227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(10), ack => type_cast_96_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_76_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_76_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_76_Sample/ra
      -- 
    ra_200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_76_inst_ack_0, ack => sendOutput_CP_26_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	58 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	47 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_76_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_76_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_76_Update/ca
      -- 
    ca_205_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_76_inst_ack_1, ack => sendOutput_CP_26_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_86_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_86_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_86_Sample/ra
      -- 
    ra_214_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_86_inst_ack_0, ack => sendOutput_CP_26_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	58 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	44 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_86_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_86_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_86_Update/ca
      -- 
    ca_219_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_86_inst_ack_1, ack => sendOutput_CP_26_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_96_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_96_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_96_Sample/ra
      -- 
    ra_228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_96_inst_ack_0, ack => sendOutput_CP_26_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	58 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	41 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_96_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_96_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_96_Update/ca
      -- 
    ca_233_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_96_inst_ack_1, ack => sendOutput_CP_26_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	10 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_106_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_106_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_106_Sample/ra
      -- 
    ra_242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_106_inst_ack_0, ack => sendOutput_CP_26_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	58 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	38 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_106_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_106_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_106_Update/ca
      -- 
    ca_247_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_106_inst_ack_1, ack => sendOutput_CP_26_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	10 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_116_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_116_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_116_Sample/ra
      -- 
    ra_256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_116_inst_ack_0, ack => sendOutput_CP_26_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	58 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	35 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_116_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_116_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_116_Update/ca
      -- 
    ca_261_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_116_inst_ack_1, ack => sendOutput_CP_26_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	10 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_126_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_126_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_126_Sample/ra
      -- 
    ra_270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_126_inst_ack_0, ack => sendOutput_CP_26_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	58 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	32 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_126_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_126_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_126_Update/ca
      -- 
    ca_275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_126_inst_ack_1, ack => sendOutput_CP_26_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	10 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_136_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_136_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_136_Sample/ra
      -- 
    ra_284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_136_inst_ack_0, ack => sendOutput_CP_26_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	58 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	29 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_136_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_136_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_136_Update/ca
      -- 
    ca_289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_136_inst_ack_1, ack => sendOutput_CP_26_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	10 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_146_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_146_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_146_Sample/ra
      -- 
    ra_298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_146_inst_ack_0, ack => sendOutput_CP_26_elements(25)); -- 
    -- CP-element group 26:  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	58 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (6) 
      -- CP-element group 26: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_146_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_146_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_146_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_148_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_148_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_148_Sample/req
      -- 
    ca_303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_146_inst_ack_1, ack => sendOutput_CP_26_elements(26)); -- 
    req_311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(26), ack => WPIPE_zeropad_output_pipe_148_inst_req_0); -- 
    -- CP-element group 27:  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (6) 
      -- CP-element group 27: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_148_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_148_update_start_
      -- CP-element group 27: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_148_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_148_Sample/ack
      -- CP-element group 27: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_148_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_148_Update/req
      -- 
    ack_312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_148_inst_ack_0, ack => sendOutput_CP_26_elements(27)); -- 
    req_316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(27), ack => WPIPE_zeropad_output_pipe_148_inst_req_1); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_148_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_148_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_148_Update/ack
      -- 
    ack_317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_148_inst_ack_1, ack => sendOutput_CP_26_elements(28)); -- 
    -- CP-element group 29:  join  transition  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: 	24 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_151_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_151_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_151_Sample/req
      -- 
    req_325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(29), ack => WPIPE_zeropad_output_pipe_151_inst_req_0); -- 
    sendOutput_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(28) & sendOutput_CP_26_elements(24);
      gj_sendOutput_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_151_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_151_update_start_
      -- CP-element group 30: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_151_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_151_Sample/ack
      -- CP-element group 30: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_151_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_151_Update/req
      -- 
    ack_326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_151_inst_ack_0, ack => sendOutput_CP_26_elements(30)); -- 
    req_330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(30), ack => WPIPE_zeropad_output_pipe_151_inst_req_1); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_151_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_151_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_151_Update/ack
      -- 
    ack_331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_151_inst_ack_1, ack => sendOutput_CP_26_elements(31)); -- 
    -- CP-element group 32:  join  transition  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: 	22 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_154_sample_start_
      -- CP-element group 32: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_154_Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_154_Sample/req
      -- 
    req_339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(32), ack => WPIPE_zeropad_output_pipe_154_inst_req_0); -- 
    sendOutput_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(31) & sendOutput_CP_26_elements(22);
      gj_sendOutput_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_154_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_154_update_start_
      -- CP-element group 33: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_154_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_154_Sample/ack
      -- CP-element group 33: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_154_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_154_Update/req
      -- 
    ack_340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_154_inst_ack_0, ack => sendOutput_CP_26_elements(33)); -- 
    req_344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(33), ack => WPIPE_zeropad_output_pipe_154_inst_req_1); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_154_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_154_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_154_Update/ack
      -- 
    ack_345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_154_inst_ack_1, ack => sendOutput_CP_26_elements(34)); -- 
    -- CP-element group 35:  join  transition  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: 	20 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_157_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_157_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_157_Sample/req
      -- 
    req_353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(35), ack => WPIPE_zeropad_output_pipe_157_inst_req_0); -- 
    sendOutput_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(34) & sendOutput_CP_26_elements(20);
      gj_sendOutput_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  transition  input  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (6) 
      -- CP-element group 36: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_157_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_157_update_start_
      -- CP-element group 36: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_157_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_157_Sample/ack
      -- CP-element group 36: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_157_Update/$entry
      -- CP-element group 36: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_157_Update/req
      -- 
    ack_354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_157_inst_ack_0, ack => sendOutput_CP_26_elements(36)); -- 
    req_358_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_358_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(36), ack => WPIPE_zeropad_output_pipe_157_inst_req_1); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_157_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_157_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_157_Update/ack
      -- 
    ack_359_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_157_inst_ack_1, ack => sendOutput_CP_26_elements(37)); -- 
    -- CP-element group 38:  join  transition  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: 	18 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_160_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_160_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_160_Sample/req
      -- 
    req_367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(38), ack => WPIPE_zeropad_output_pipe_160_inst_req_0); -- 
    sendOutput_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(37) & sendOutput_CP_26_elements(18);
      gj_sendOutput_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (6) 
      -- CP-element group 39: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_160_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_160_update_start_
      -- CP-element group 39: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_160_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_160_Sample/ack
      -- CP-element group 39: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_160_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_160_Update/req
      -- 
    ack_368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_160_inst_ack_0, ack => sendOutput_CP_26_elements(39)); -- 
    req_372_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_372_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(39), ack => WPIPE_zeropad_output_pipe_160_inst_req_1); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_160_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_160_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_160_Update/ack
      -- 
    ack_373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_160_inst_ack_1, ack => sendOutput_CP_26_elements(40)); -- 
    -- CP-element group 41:  join  transition  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: 	16 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_163_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_163_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_163_Sample/req
      -- 
    req_381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(41), ack => WPIPE_zeropad_output_pipe_163_inst_req_0); -- 
    sendOutput_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(40) & sendOutput_CP_26_elements(16);
      gj_sendOutput_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (6) 
      -- CP-element group 42: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_163_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_163_update_start_
      -- CP-element group 42: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_163_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_163_Sample/ack
      -- CP-element group 42: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_163_Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_163_Update/req
      -- 
    ack_382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_163_inst_ack_0, ack => sendOutput_CP_26_elements(42)); -- 
    req_386_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_386_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(42), ack => WPIPE_zeropad_output_pipe_163_inst_req_1); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_163_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_163_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_163_Update/ack
      -- 
    ack_387_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_163_inst_ack_1, ack => sendOutput_CP_26_elements(43)); -- 
    -- CP-element group 44:  join  transition  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: 	14 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_166_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_166_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_166_Sample/req
      -- 
    req_395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(44), ack => WPIPE_zeropad_output_pipe_166_inst_req_0); -- 
    sendOutput_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(43) & sendOutput_CP_26_elements(14);
      gj_sendOutput_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_166_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_166_update_start_
      -- CP-element group 45: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_166_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_166_Sample/ack
      -- CP-element group 45: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_166_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_166_Update/req
      -- 
    ack_396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_166_inst_ack_0, ack => sendOutput_CP_26_elements(45)); -- 
    req_400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(45), ack => WPIPE_zeropad_output_pipe_166_inst_req_1); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_166_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_166_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_166_Update/ack
      -- 
    ack_401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_166_inst_ack_1, ack => sendOutput_CP_26_elements(46)); -- 
    -- CP-element group 47:  join  transition  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: 	12 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_169_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_169_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_169_Sample/req
      -- 
    req_409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(47), ack => WPIPE_zeropad_output_pipe_169_inst_req_0); -- 
    sendOutput_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(46) & sendOutput_CP_26_elements(12);
      gj_sendOutput_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (6) 
      -- CP-element group 48: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_169_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_169_update_start_
      -- CP-element group 48: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_169_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_169_Sample/ack
      -- CP-element group 48: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_169_Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_169_Update/req
      -- 
    ack_410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_169_inst_ack_0, ack => sendOutput_CP_26_elements(48)); -- 
    req_414_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_414_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(48), ack => WPIPE_zeropad_output_pipe_169_inst_req_1); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_169_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_169_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/WPIPE_zeropad_output_pipe_169_Update/ack
      -- 
    ack_415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_169_inst_ack_1, ack => sendOutput_CP_26_elements(49)); -- 
    -- CP-element group 50:  branch  join  transition  place  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: 	5 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (10) 
      -- CP-element group 50: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182__exit__
      -- CP-element group 50: 	 branch_block_stmt_22/if_stmt_183__entry__
      -- CP-element group 50: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/$exit
      -- CP-element group 50: 	 branch_block_stmt_22/if_stmt_183_dead_link/$entry
      -- CP-element group 50: 	 branch_block_stmt_22/if_stmt_183_eval_test/$entry
      -- CP-element group 50: 	 branch_block_stmt_22/if_stmt_183_eval_test/$exit
      -- CP-element group 50: 	 branch_block_stmt_22/if_stmt_183_eval_test/branch_req
      -- CP-element group 50: 	 branch_block_stmt_22/R_exitcond2_184_place
      -- CP-element group 50: 	 branch_block_stmt_22/if_stmt_183_if_link/$entry
      -- CP-element group 50: 	 branch_block_stmt_22/if_stmt_183_else_link/$entry
      -- 
    branch_req_423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(50), ack => if_stmt_183_branch_req_0); -- 
    sendOutput_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(49) & sendOutput_CP_26_elements(5);
      gj_sendOutput_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  merge  transition  place  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	59 
    -- CP-element group 51:  members (13) 
      -- CP-element group 51: 	 branch_block_stmt_22/merge_stmt_189__exit__
      -- CP-element group 51: 	 branch_block_stmt_22/forx_xendx_xloopexit_forx_xend
      -- CP-element group 51: 	 branch_block_stmt_22/if_stmt_183_if_link/$exit
      -- CP-element group 51: 	 branch_block_stmt_22/if_stmt_183_if_link/if_choice_transition
      -- CP-element group 51: 	 branch_block_stmt_22/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 51: 	 branch_block_stmt_22/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 51: 	 branch_block_stmt_22/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 51: 	 branch_block_stmt_22/merge_stmt_189_PhiReqMerge
      -- CP-element group 51: 	 branch_block_stmt_22/merge_stmt_189_PhiAck/$entry
      -- CP-element group 51: 	 branch_block_stmt_22/merge_stmt_189_PhiAck/$exit
      -- CP-element group 51: 	 branch_block_stmt_22/merge_stmt_189_PhiAck/dummy
      -- CP-element group 51: 	 branch_block_stmt_22/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 51: 	 branch_block_stmt_22/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_183_branch_ack_1, ack => sendOutput_CP_26_elements(51)); -- 
    -- CP-element group 52:  fork  transition  place  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52: 	55 
    -- CP-element group 52:  members (12) 
      -- CP-element group 52: 	 branch_block_stmt_22/if_stmt_183_else_link/$exit
      -- CP-element group 52: 	 branch_block_stmt_22/if_stmt_183_else_link/else_choice_transition
      -- CP-element group 52: 	 branch_block_stmt_22/forx_xbody_forx_xbody
      -- CP-element group 52: 	 branch_block_stmt_22/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 52: 	 branch_block_stmt_22/forx_xbody_forx_xbody_PhiReq/phi_stmt_55/$entry
      -- CP-element group 52: 	 branch_block_stmt_22/forx_xbody_forx_xbody_PhiReq/phi_stmt_55/phi_stmt_55_sources/$entry
      -- CP-element group 52: 	 branch_block_stmt_22/forx_xbody_forx_xbody_PhiReq/phi_stmt_55/phi_stmt_55_sources/type_cast_58/$entry
      -- CP-element group 52: 	 branch_block_stmt_22/forx_xbody_forx_xbody_PhiReq/phi_stmt_55/phi_stmt_55_sources/type_cast_58/SplitProtocol/$entry
      -- CP-element group 52: 	 branch_block_stmt_22/forx_xbody_forx_xbody_PhiReq/phi_stmt_55/phi_stmt_55_sources/type_cast_58/SplitProtocol/Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_22/forx_xbody_forx_xbody_PhiReq/phi_stmt_55/phi_stmt_55_sources/type_cast_58/SplitProtocol/Sample/rr
      -- CP-element group 52: 	 branch_block_stmt_22/forx_xbody_forx_xbody_PhiReq/phi_stmt_55/phi_stmt_55_sources/type_cast_58/SplitProtocol/Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_22/forx_xbody_forx_xbody_PhiReq/phi_stmt_55/phi_stmt_55_sources/type_cast_58/SplitProtocol/Update/cr
      -- 
    else_choice_transition_432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_183_branch_ack_0, ack => sendOutput_CP_26_elements(52)); -- 
    rr_476_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_476_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(52), ack => type_cast_58_inst_req_0); -- 
    cr_481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(52), ack => type_cast_58_inst_req_1); -- 
    -- CP-element group 53:  transition  output  delay-element  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	4 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	57 
    -- CP-element group 53:  members (5) 
      -- CP-element group 53: 	 branch_block_stmt_22/bbx_xnph_forx_xbody_PhiReq/$exit
      -- CP-element group 53: 	 branch_block_stmt_22/bbx_xnph_forx_xbody_PhiReq/phi_stmt_55/$exit
      -- CP-element group 53: 	 branch_block_stmt_22/bbx_xnph_forx_xbody_PhiReq/phi_stmt_55/phi_stmt_55_sources/$exit
      -- CP-element group 53: 	 branch_block_stmt_22/bbx_xnph_forx_xbody_PhiReq/phi_stmt_55/phi_stmt_55_sources/type_cast_61_konst_delay_trans
      -- CP-element group 53: 	 branch_block_stmt_22/bbx_xnph_forx_xbody_PhiReq/phi_stmt_55/phi_stmt_55_req
      -- 
    phi_stmt_55_req_457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_55_req_457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(53), ack => phi_stmt_55_req_1); -- 
    -- Element group sendOutput_CP_26_elements(53) is a control-delay.
    cp_element_53_delay: control_delay_element  generic map(name => " 53_delay", delay_value => 1)  port map(req => sendOutput_CP_26_elements(4), ack => sendOutput_CP_26_elements(53), clk => clk, reset =>reset);
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (2) 
      -- CP-element group 54: 	 branch_block_stmt_22/forx_xbody_forx_xbody_PhiReq/phi_stmt_55/phi_stmt_55_sources/type_cast_58/SplitProtocol/Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_22/forx_xbody_forx_xbody_PhiReq/phi_stmt_55/phi_stmt_55_sources/type_cast_58/SplitProtocol/Sample/ra
      -- 
    ra_477_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_58_inst_ack_0, ack => sendOutput_CP_26_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	52 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (2) 
      -- CP-element group 55: 	 branch_block_stmt_22/forx_xbody_forx_xbody_PhiReq/phi_stmt_55/phi_stmt_55_sources/type_cast_58/SplitProtocol/Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_22/forx_xbody_forx_xbody_PhiReq/phi_stmt_55/phi_stmt_55_sources/type_cast_58/SplitProtocol/Update/ca
      -- 
    ca_482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_58_inst_ack_1, ack => sendOutput_CP_26_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (6) 
      -- CP-element group 56: 	 branch_block_stmt_22/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 56: 	 branch_block_stmt_22/forx_xbody_forx_xbody_PhiReq/phi_stmt_55/$exit
      -- CP-element group 56: 	 branch_block_stmt_22/forx_xbody_forx_xbody_PhiReq/phi_stmt_55/phi_stmt_55_sources/$exit
      -- CP-element group 56: 	 branch_block_stmt_22/forx_xbody_forx_xbody_PhiReq/phi_stmt_55/phi_stmt_55_sources/type_cast_58/$exit
      -- CP-element group 56: 	 branch_block_stmt_22/forx_xbody_forx_xbody_PhiReq/phi_stmt_55/phi_stmt_55_sources/type_cast_58/SplitProtocol/$exit
      -- CP-element group 56: 	 branch_block_stmt_22/forx_xbody_forx_xbody_PhiReq/phi_stmt_55/phi_stmt_55_req
      -- 
    phi_stmt_55_req_483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_55_req_483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(56), ack => phi_stmt_55_req_0); -- 
    sendOutput_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(54) & sendOutput_CP_26_elements(55);
      gj_sendOutput_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  merge  transition  place  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	53 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (2) 
      -- CP-element group 57: 	 branch_block_stmt_22/merge_stmt_54_PhiReqMerge
      -- CP-element group 57: 	 branch_block_stmt_22/merge_stmt_54_PhiAck/$entry
      -- 
    sendOutput_CP_26_elements(57) <= OrReduce(sendOutput_CP_26_elements(53) & sendOutput_CP_26_elements(56));
    -- CP-element group 58:  fork  transition  place  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	16 
    -- CP-element group 58: 	5 
    -- CP-element group 58: 	14 
    -- CP-element group 58: 	6 
    -- CP-element group 58: 	22 
    -- CP-element group 58: 	18 
    -- CP-element group 58: 	10 
    -- CP-element group 58: 	12 
    -- CP-element group 58: 	8 
    -- CP-element group 58: 	26 
    -- CP-element group 58: 	20 
    -- CP-element group 58: 	24 
    -- CP-element group 58:  members (53) 
      -- CP-element group 58: 	 branch_block_stmt_22/merge_stmt_54__exit__
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182__entry__
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_76_update_start_
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/$entry
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/addr_of_68_update_start_
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/array_obj_ref_67_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/array_obj_ref_67_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/array_obj_ref_67_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/array_obj_ref_67_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/array_obj_ref_67_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/array_obj_ref_67_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/array_obj_ref_67_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/array_obj_ref_67_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/array_obj_ref_67_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/array_obj_ref_67_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/array_obj_ref_67_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/array_obj_ref_67_final_index_sum_regn_update_start
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/array_obj_ref_67_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/array_obj_ref_67_final_index_sum_regn_Sample/req
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/array_obj_ref_67_final_index_sum_regn_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/array_obj_ref_67_final_index_sum_regn_Update/req
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/addr_of_68_complete/$entry
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/addr_of_68_complete/req
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/ptr_deref_72_update_start_
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/ptr_deref_72_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/ptr_deref_72_Update/word_access_complete/$entry
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/ptr_deref_72_Update/word_access_complete/word_0/$entry
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/ptr_deref_72_Update/word_access_complete/word_0/cr
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_76_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_76_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_86_update_start_
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_86_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_86_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_96_update_start_
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_96_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_96_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_106_update_start_
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_106_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_106_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_116_update_start_
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_116_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_116_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_126_update_start_
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_126_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_126_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_136_update_start_
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_136_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_136_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_146_update_start_
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_146_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_22/assign_stmt_69_to_assign_stmt_182/type_cast_146_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_22/merge_stmt_54_PhiAck/$exit
      -- CP-element group 58: 	 branch_block_stmt_22/merge_stmt_54_PhiAck/phi_stmt_55_ack
      -- 
    phi_stmt_55_ack_488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_55_ack_0, ack => sendOutput_CP_26_elements(58)); -- 
    req_120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => array_obj_ref_67_index_offset_req_0); -- 
    req_125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => array_obj_ref_67_index_offset_req_1); -- 
    req_140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => addr_of_68_final_reg_req_1); -- 
    cr_185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => ptr_deref_72_load_0_req_1); -- 
    cr_204_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_204_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => type_cast_76_inst_req_1); -- 
    cr_218_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_218_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => type_cast_86_inst_req_1); -- 
    cr_232_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_232_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => type_cast_96_inst_req_1); -- 
    cr_246_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_246_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => type_cast_106_inst_req_1); -- 
    cr_260_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_260_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => type_cast_116_inst_req_1); -- 
    cr_274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => type_cast_126_inst_req_1); -- 
    cr_288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => type_cast_136_inst_req_1); -- 
    cr_302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => type_cast_146_inst_req_1); -- 
    -- CP-element group 59:  merge  transition  place  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	51 
    -- CP-element group 59: 	2 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (16) 
      -- CP-element group 59: 	 $exit
      -- CP-element group 59: 	 branch_block_stmt_22/$exit
      -- CP-element group 59: 	 branch_block_stmt_22/branch_block_stmt_22__exit__
      -- CP-element group 59: 	 branch_block_stmt_22/merge_stmt_191__exit__
      -- CP-element group 59: 	 branch_block_stmt_22/return__
      -- CP-element group 59: 	 branch_block_stmt_22/merge_stmt_193__exit__
      -- CP-element group 59: 	 branch_block_stmt_22/merge_stmt_191_PhiReqMerge
      -- CP-element group 59: 	 branch_block_stmt_22/merge_stmt_191_PhiAck/$entry
      -- CP-element group 59: 	 branch_block_stmt_22/merge_stmt_191_PhiAck/$exit
      -- CP-element group 59: 	 branch_block_stmt_22/merge_stmt_191_PhiAck/dummy
      -- CP-element group 59: 	 branch_block_stmt_22/return___PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_22/return___PhiReq/$exit
      -- CP-element group 59: 	 branch_block_stmt_22/merge_stmt_193_PhiReqMerge
      -- CP-element group 59: 	 branch_block_stmt_22/merge_stmt_193_PhiAck/$entry
      -- CP-element group 59: 	 branch_block_stmt_22/merge_stmt_193_PhiAck/$exit
      -- CP-element group 59: 	 branch_block_stmt_22/merge_stmt_193_PhiAck/dummy
      -- 
    sendOutput_CP_26_elements(59) <= OrReduce(sendOutput_CP_26_elements(51) & sendOutput_CP_26_elements(2));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_30_wire : std_logic_vector(31 downto 0);
    signal R_indvar_66_resized : std_logic_vector(13 downto 0);
    signal R_indvar_66_scaled : std_logic_vector(13 downto 0);
    signal array_obj_ref_67_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_67_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_67_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_67_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_67_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_67_root_address : std_logic_vector(13 downto 0);
    signal arrayidx_69 : std_logic_vector(31 downto 0);
    signal cmp68_41 : std_logic_vector(0 downto 0);
    signal conv12_87 : std_logic_vector(7 downto 0);
    signal conv18_97 : std_logic_vector(7 downto 0);
    signal conv24_107 : std_logic_vector(7 downto 0);
    signal conv30_117 : std_logic_vector(7 downto 0);
    signal conv36_127 : std_logic_vector(7 downto 0);
    signal conv42_137 : std_logic_vector(7 downto 0);
    signal conv48_147 : std_logic_vector(7 downto 0);
    signal conv_77 : std_logic_vector(7 downto 0);
    signal exitcond2_182 : std_logic_vector(0 downto 0);
    signal indvar_55 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_177 : std_logic_vector(63 downto 0);
    signal ptr_deref_72_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_72_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_72_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_72_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_72_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr15_93 : std_logic_vector(63 downto 0);
    signal shr21_103 : std_logic_vector(63 downto 0);
    signal shr27_113 : std_logic_vector(63 downto 0);
    signal shr33_123 : std_logic_vector(63 downto 0);
    signal shr39_133 : std_logic_vector(63 downto 0);
    signal shr45_143 : std_logic_vector(63 downto 0);
    signal shr67_32 : std_logic_vector(31 downto 0);
    signal shr9_83 : std_logic_vector(63 downto 0);
    signal tmp1_52 : std_logic_vector(63 downto 0);
    signal tmp4_73 : std_logic_vector(63 downto 0);
    signal type_cast_101_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_111_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_121_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_131_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_141_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_175_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_26_wire : std_logic_vector(31 downto 0);
    signal type_cast_29_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_35_wire : std_logic_vector(31 downto 0);
    signal type_cast_38_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_58_wire : std_logic_vector(63 downto 0);
    signal type_cast_61_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_81_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_91_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_67_constant_part_of_offset <= "00000000000000";
    array_obj_ref_67_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_67_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_67_resized_base_address <= "00000000000000";
    ptr_deref_72_word_offset_0 <= "00000000000000";
    type_cast_101_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_111_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_121_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_131_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_141_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_175_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_29_wire_constant <= "00000000000000000000000000000010";
    type_cast_38_wire_constant <= "00000000000000000000000000000000";
    type_cast_61_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_81_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_91_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    phi_stmt_55: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_58_wire & type_cast_61_wire_constant;
      req <= phi_stmt_55_req_0 & phi_stmt_55_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_55",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_55_ack_0,
          idata => idata,
          odata => indvar_55,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_55
    addr_of_68_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_68_final_reg_req_0;
      addr_of_68_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_68_final_reg_req_1;
      addr_of_68_final_reg_ack_1<= rack(0);
      addr_of_68_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_68_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_67_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_69,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_106_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_106_inst_req_0;
      type_cast_106_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_106_inst_req_1;
      type_cast_106_inst_ack_1<= rack(0);
      type_cast_106_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_106_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr21_103,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv24_107,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_116_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_116_inst_req_0;
      type_cast_116_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_116_inst_req_1;
      type_cast_116_inst_ack_1<= rack(0);
      type_cast_116_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_116_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr27_113,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv30_117,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_126_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_126_inst_req_0;
      type_cast_126_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_126_inst_req_1;
      type_cast_126_inst_ack_1<= rack(0);
      type_cast_126_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_126_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr33_123,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv36_127,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_136_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_136_inst_req_0;
      type_cast_136_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_136_inst_req_1;
      type_cast_136_inst_ack_1<= rack(0);
      type_cast_136_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_136_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr39_133,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv42_137,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_146_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_146_inst_req_0;
      type_cast_146_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_146_inst_req_1;
      type_cast_146_inst_ack_1<= rack(0);
      type_cast_146_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_146_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr45_143,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv48_147,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_26_inst
    process(size_buffer) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := size_buffer(31 downto 0);
      type_cast_26_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_31_inst
    process(ASHR_i32_i32_30_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_30_wire(31 downto 0);
      shr67_32 <= tmp_var; -- 
    end process;
    -- interlock type_cast_35_inst
    process(shr67_32) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := shr67_32(31 downto 0);
      type_cast_35_wire <= tmp_var; -- 
    end process;
    type_cast_51_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_51_inst_req_0;
      type_cast_51_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_51_inst_req_1;
      type_cast_51_inst_ack_1<= rack(0);
      type_cast_51_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_51_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr67_32,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp1_52,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_58_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_58_inst_req_0;
      type_cast_58_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_58_inst_req_1;
      type_cast_58_inst_ack_1<= rack(0);
      type_cast_58_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_58_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_177,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_58_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_76_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_76_inst_req_0;
      type_cast_76_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_76_inst_req_1;
      type_cast_76_inst_ack_1<= rack(0);
      type_cast_76_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_76_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp4_73,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_77,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_86_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_86_inst_req_0;
      type_cast_86_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_86_inst_req_1;
      type_cast_86_inst_ack_1<= rack(0);
      type_cast_86_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_86_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr9_83,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv12_87,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_96_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_96_inst_req_0;
      type_cast_96_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_96_inst_req_1;
      type_cast_96_inst_ack_1<= rack(0);
      type_cast_96_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_96_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr15_93,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv18_97,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_67_index_1_rename
    process(R_indvar_66_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_66_resized;
      ov(13 downto 0) := iv;
      R_indvar_66_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_67_index_1_resize
    process(indvar_55) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_55;
      ov := iv(13 downto 0);
      R_indvar_66_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_67_root_address_inst
    process(array_obj_ref_67_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_67_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_67_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_72_addr_0
    process(ptr_deref_72_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_72_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_72_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_72_base_resize
    process(arrayidx_69) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_69;
      ov := iv(13 downto 0);
      ptr_deref_72_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_72_gather_scatter
    process(ptr_deref_72_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_72_data_0;
      ov(63 downto 0) := iv;
      tmp4_73 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_72_root_address_inst
    process(ptr_deref_72_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_72_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_72_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_183_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond2_182;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_183_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_183_branch_req_0,
          ack0 => if_stmt_183_branch_ack_0,
          ack1 => if_stmt_183_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_42_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp68_41;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_42_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_42_branch_req_0,
          ack0 => if_stmt_42_branch_ack_0,
          ack1 => if_stmt_42_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_176_inst
    process(indvar_55) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_55, type_cast_175_wire_constant, tmp_var);
      indvarx_xnext_177 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_30_inst
    process(type_cast_26_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_26_wire, type_cast_29_wire_constant, tmp_var);
      ASHR_i32_i32_30_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_181_inst
    process(indvarx_xnext_177, tmp1_52) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_177, tmp1_52, tmp_var);
      exitcond2_182 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_102_inst
    process(tmp4_73) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_73, type_cast_101_wire_constant, tmp_var);
      shr21_103 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_112_inst
    process(tmp4_73) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_73, type_cast_111_wire_constant, tmp_var);
      shr27_113 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_122_inst
    process(tmp4_73) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_73, type_cast_121_wire_constant, tmp_var);
      shr33_123 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_132_inst
    process(tmp4_73) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_73, type_cast_131_wire_constant, tmp_var);
      shr39_133 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_142_inst
    process(tmp4_73) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_73, type_cast_141_wire_constant, tmp_var);
      shr45_143 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_82_inst
    process(tmp4_73) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_73, type_cast_81_wire_constant, tmp_var);
      shr9_83 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_92_inst
    process(tmp4_73) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_73, type_cast_91_wire_constant, tmp_var);
      shr15_93 <= tmp_var; --
    end process;
    -- binary operator SGT_i32_u1_39_inst
    process(type_cast_35_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(type_cast_35_wire, type_cast_38_wire_constant, tmp_var);
      cmp68_41 <= tmp_var; --
    end process;
    -- shared split operator group (11) : array_obj_ref_67_index_offset 
    ApIntAdd_group_11: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_66_scaled;
      array_obj_ref_67_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_67_index_offset_req_0;
      array_obj_ref_67_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_67_index_offset_req_1;
      array_obj_ref_67_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_11_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_11_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_11",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared load operator group (0) : ptr_deref_72_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_72_load_0_req_0;
      ptr_deref_72_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_72_load_0_req_1;
      ptr_deref_72_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_72_word_address_0;
      ptr_deref_72_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared outport operator group (0) : WPIPE_zeropad_output_pipe_148_inst WPIPE_zeropad_output_pipe_151_inst WPIPE_zeropad_output_pipe_154_inst WPIPE_zeropad_output_pipe_157_inst WPIPE_zeropad_output_pipe_160_inst WPIPE_zeropad_output_pipe_163_inst WPIPE_zeropad_output_pipe_166_inst WPIPE_zeropad_output_pipe_169_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 7 downto 0);
      signal update_req, update_ack : BooleanArray( 7 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 7 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      sample_req_unguarded(7) <= WPIPE_zeropad_output_pipe_148_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_zeropad_output_pipe_151_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_zeropad_output_pipe_154_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_zeropad_output_pipe_157_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_zeropad_output_pipe_160_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_zeropad_output_pipe_163_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_zeropad_output_pipe_166_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_zeropad_output_pipe_169_inst_req_0;
      WPIPE_zeropad_output_pipe_148_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_zeropad_output_pipe_151_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_zeropad_output_pipe_154_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_zeropad_output_pipe_157_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_zeropad_output_pipe_160_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_zeropad_output_pipe_163_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_zeropad_output_pipe_166_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_zeropad_output_pipe_169_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(7) <= WPIPE_zeropad_output_pipe_148_inst_req_1;
      update_req_unguarded(6) <= WPIPE_zeropad_output_pipe_151_inst_req_1;
      update_req_unguarded(5) <= WPIPE_zeropad_output_pipe_154_inst_req_1;
      update_req_unguarded(4) <= WPIPE_zeropad_output_pipe_157_inst_req_1;
      update_req_unguarded(3) <= WPIPE_zeropad_output_pipe_160_inst_req_1;
      update_req_unguarded(2) <= WPIPE_zeropad_output_pipe_163_inst_req_1;
      update_req_unguarded(1) <= WPIPE_zeropad_output_pipe_166_inst_req_1;
      update_req_unguarded(0) <= WPIPE_zeropad_output_pipe_169_inst_req_1;
      WPIPE_zeropad_output_pipe_148_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_zeropad_output_pipe_151_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_zeropad_output_pipe_154_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_zeropad_output_pipe_157_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_zeropad_output_pipe_160_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_zeropad_output_pipe_163_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_zeropad_output_pipe_166_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_zeropad_output_pipe_169_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      data_in <= conv48_147 & conv42_137 & conv36_127 & conv30_117 & conv24_107 & conv18_97 & conv12_87 & conv_77;
      zeropad_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "zeropad_output_pipe_write_0_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      zeropad_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "zeropad_output_pipe", data_width => 8, num_reqs => 8, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => zeropad_output_pipe_pipe_write_req(0),
          oack => zeropad_output_pipe_pipe_write_ack(0),
          odata => zeropad_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end sendOutput_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    c : out  std_logic_vector(63 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal c_buffer :  std_logic_vector(63 downto 0);
  signal c_update_enable: Boolean;
  signal timer_CP_520_start: Boolean;
  signal timer_CP_520_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal LOAD_count_199_load_0_req_0 : boolean;
  signal LOAD_count_199_load_0_ack_0 : boolean;
  signal LOAD_count_199_load_0_req_1 : boolean;
  signal LOAD_count_199_load_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_520_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= c_buffer;
  c <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_520_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_520_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_520_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_520: Block -- control-path 
    signal timer_CP_520_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    timer_CP_520_elements(0) <= timer_CP_520_start;
    timer_CP_520_symbol <= timer_CP_520_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_200/$entry
      -- CP-element group 0: 	 assign_stmt_200/LOAD_count_199_sample_start_
      -- CP-element group 0: 	 assign_stmt_200/LOAD_count_199_update_start_
      -- CP-element group 0: 	 assign_stmt_200/LOAD_count_199_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_200/LOAD_count_199_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_200/LOAD_count_199_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_200/LOAD_count_199_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_200/LOAD_count_199_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_200/LOAD_count_199_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_200/LOAD_count_199_Update/$entry
      -- CP-element group 0: 	 assign_stmt_200/LOAD_count_199_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_200/LOAD_count_199_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_200/LOAD_count_199_Update/word_access_complete/word_0/cr
      -- 
    cr_552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_520_elements(0), ack => LOAD_count_199_load_0_req_1); -- 
    rr_541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_520_elements(0), ack => LOAD_count_199_load_0_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 assign_stmt_200/LOAD_count_199_sample_completed_
      -- CP-element group 1: 	 assign_stmt_200/LOAD_count_199_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_200/LOAD_count_199_Sample/word_access_start/$exit
      -- CP-element group 1: 	 assign_stmt_200/LOAD_count_199_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 assign_stmt_200/LOAD_count_199_Sample/word_access_start/word_0/ra
      -- 
    ra_542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_199_load_0_ack_0, ack => timer_CP_520_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_200/$exit
      -- CP-element group 2: 	 assign_stmt_200/LOAD_count_199_update_completed_
      -- CP-element group 2: 	 assign_stmt_200/LOAD_count_199_Update/$exit
      -- CP-element group 2: 	 assign_stmt_200/LOAD_count_199_Update/word_access_complete/$exit
      -- CP-element group 2: 	 assign_stmt_200/LOAD_count_199_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 assign_stmt_200/LOAD_count_199_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 assign_stmt_200/LOAD_count_199_Update/LOAD_count_199_Merge/$entry
      -- CP-element group 2: 	 assign_stmt_200/LOAD_count_199_Update/LOAD_count_199_Merge/$exit
      -- CP-element group 2: 	 assign_stmt_200/LOAD_count_199_Update/LOAD_count_199_Merge/merge_req
      -- CP-element group 2: 	 assign_stmt_200/LOAD_count_199_Update/LOAD_count_199_Merge/merge_ack
      -- 
    ca_553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_199_load_0_ack_1, ack => timer_CP_520_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_count_199_data_0 : std_logic_vector(63 downto 0);
    signal LOAD_count_199_word_address_0 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    LOAD_count_199_word_address_0 <= "0";
    -- equivalence LOAD_count_199_gather_scatter
    process(LOAD_count_199_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_count_199_data_0;
      ov(63 downto 0) := iv;
      c_buffer <= ov(63 downto 0);
      --
    end process;
    -- shared load operator group (0) : LOAD_count_199_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_count_199_load_0_req_0;
      LOAD_count_199_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_count_199_load_0_req_1;
      LOAD_count_199_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_count_199_word_address_0;
      LOAD_count_199_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(0 downto 0),
          mtag => memory_space_2_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(63 downto 0),
          mtag => memory_space_2_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timerDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timerDaemon;
architecture timerDaemon_arch of timerDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal timerDaemon_CP_559_start: Boolean;
  signal timerDaemon_CP_559_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal do_while_stmt_204_branch_req_0 : boolean;
  signal STORE_count_214_store_0_req_1 : boolean;
  signal STORE_count_214_store_0_ack_1 : boolean;
  signal phi_stmt_206_ack_0 : boolean;
  signal do_while_stmt_204_branch_ack_0 : boolean;
  signal ADD_u64_u64_210_inst_ack_1 : boolean;
  signal STORE_count_214_store_0_ack_0 : boolean;
  signal ADD_u64_u64_210_inst_req_1 : boolean;
  signal STORE_count_214_store_0_req_0 : boolean;
  signal ADD_u64_u64_210_inst_ack_0 : boolean;
  signal ADD_u64_u64_210_inst_req_0 : boolean;
  signal phi_stmt_206_req_1 : boolean;
  signal phi_stmt_206_req_0 : boolean;
  signal do_while_stmt_204_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timerDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timerDaemon_CP_559_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timerDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_559_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timerDaemon_CP_559_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_559_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timerDaemon_CP_559: Block -- control-path 
    signal timerDaemon_CP_559_elements: BooleanArray(39 downto 0);
    -- 
  begin -- 
    timerDaemon_CP_559_elements(0) <= timerDaemon_CP_559_start;
    timerDaemon_CP_559_symbol <= timerDaemon_CP_559_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_203/do_while_stmt_204__entry__
      -- CP-element group 0: 	 branch_block_stmt_203/branch_block_stmt_203__entry__
      -- CP-element group 0: 	 branch_block_stmt_203/$entry
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	39 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_203/do_while_stmt_204__exit__
      -- CP-element group 1: 	 branch_block_stmt_203/branch_block_stmt_203__exit__
      -- CP-element group 1: 	 branch_block_stmt_203/$exit
      -- CP-element group 1: 	 $exit
      -- 
    timerDaemon_CP_559_elements(1) <= timerDaemon_CP_559_elements(39);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204__entry__
      -- CP-element group 2: 	 branch_block_stmt_203/do_while_stmt_204/$entry
      -- 
    timerDaemon_CP_559_elements(2) <= timerDaemon_CP_559_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	39 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204__exit__
      -- 
    -- Element group timerDaemon_CP_559_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_203/do_while_stmt_204/loop_back
      -- 
    -- Element group timerDaemon_CP_559_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	37 
    -- CP-element group 5: 	38 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_203/do_while_stmt_204/condition_done
      -- CP-element group 5: 	 branch_block_stmt_203/do_while_stmt_204/loop_taken/$entry
      -- CP-element group 5: 	 branch_block_stmt_203/do_while_stmt_204/loop_exit/$entry
      -- 
    timerDaemon_CP_559_elements(5) <= timerDaemon_CP_559_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	36 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_203/do_while_stmt_204/loop_body_done
      -- 
    timerDaemon_CP_559_elements(6) <= timerDaemon_CP_559_elements(36);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	16 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/back_edge_to_loop_body
      -- 
    timerDaemon_CP_559_elements(7) <= timerDaemon_CP_559_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	18 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/first_time_through_loop_body
      -- 
    timerDaemon_CP_559_elements(8) <= timerDaemon_CP_559_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	12 
    -- CP-element group 9: 	13 
    -- CP-element group 9: 	31 
    -- CP-element group 9: 	35 
    -- CP-element group 9:  members (4) 
      -- CP-element group 9: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/STORE_count_214_root_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/STORE_count_214_word_address_calculated
      -- 
    -- Element group timerDaemon_CP_559_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: 	35 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/condition_evaluated
      -- 
    condition_evaluated_583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_559_elements(10), ack => do_while_stmt_204_branch_req_0); -- 
    timerDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 3);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_559_elements(15) & timerDaemon_CP_559_elements(35);
      gj_timerDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_559_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/phi_stmt_206_sample_start__ps
      -- CP-element group 11: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/aggregated_phi_sample_req
      -- 
    timerDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_559_elements(12) & timerDaemon_CP_559_elements(15);
      gj_timerDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_559_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: marked-predecessors 
    -- CP-element group 12: 	14 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	11 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/phi_stmt_206_sample_start_
      -- 
    timerDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_559_elements(9) & timerDaemon_CP_559_elements(14);
      gj_timerDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_559_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	9 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	33 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/phi_stmt_206_update_start__ps
      -- CP-element group 13: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/phi_stmt_206_update_start_
      -- CP-element group 13: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/aggregated_phi_update_req
      -- 
    timerDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_559_elements(9) & timerDaemon_CP_559_elements(33);
      gj_timerDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_559_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	36 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	12 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/phi_stmt_206_sample_completed__ps
      -- CP-element group 14: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/phi_stmt_206_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/aggregated_phi_sample_ack
      -- 
    -- Element group timerDaemon_CP_559_elements(14) is bound as output of CP function.
    -- CP-element group 15:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: 	31 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/phi_stmt_206_update_completed__ps
      -- CP-element group 15: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/phi_stmt_206_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/aggregated_phi_update_ack
      -- 
    -- Element group timerDaemon_CP_559_elements(15) is bound as output of CP function.
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	7 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/phi_stmt_206_loopback_trigger
      -- 
    timerDaemon_CP_559_elements(16) <= timerDaemon_CP_559_elements(7);
    -- CP-element group 17:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/phi_stmt_206_loopback_sample_req_ps
      -- CP-element group 17: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/phi_stmt_206_loopback_sample_req
      -- 
    phi_stmt_206_loopback_sample_req_598_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_206_loopback_sample_req_598_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_559_elements(17), ack => phi_stmt_206_req_0); -- 
    -- Element group timerDaemon_CP_559_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	8 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/phi_stmt_206_entry_trigger
      -- 
    timerDaemon_CP_559_elements(18) <= timerDaemon_CP_559_elements(8);
    -- CP-element group 19:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/phi_stmt_206_entry_sample_req_ps
      -- CP-element group 19: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/phi_stmt_206_entry_sample_req
      -- 
    phi_stmt_206_entry_sample_req_601_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_206_entry_sample_req_601_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_559_elements(19), ack => phi_stmt_206_req_1); -- 
    -- Element group timerDaemon_CP_559_elements(19) is bound as output of CP function.
    -- CP-element group 20:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/phi_stmt_206_phi_mux_ack
      -- CP-element group 20: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/phi_stmt_206_phi_mux_ack_ps
      -- 
    phi_stmt_206_phi_mux_ack_604_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_206_ack_0, ack => timerDaemon_CP_559_elements(20)); -- 
    -- CP-element group 21:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	23 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/ADD_u64_u64_210_sample_start__ps
      -- 
    -- Element group timerDaemon_CP_559_elements(21) is bound as output of CP function.
    -- CP-element group 22:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/ADD_u64_u64_210_update_start__ps
      -- 
    -- Element group timerDaemon_CP_559_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	21 
    -- CP-element group 23: marked-predecessors 
    -- CP-element group 23: 	25 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	25 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/ADD_u64_u64_210_Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/ADD_u64_u64_210_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/ADD_u64_u64_210_sample_start_
      -- 
    rr_617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_559_elements(23), ack => ADD_u64_u64_210_inst_req_0); -- 
    timerDaemon_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_559_elements(21) & timerDaemon_CP_559_elements(25);
      gj_timerDaemon_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_559_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	26 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/ADD_u64_u64_210_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/ADD_u64_u64_210_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/ADD_u64_u64_210_update_start_
      -- 
    cr_622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_559_elements(24), ack => ADD_u64_u64_210_inst_req_1); -- 
    timerDaemon_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_559_elements(22) & timerDaemon_CP_559_elements(26);
      gj_timerDaemon_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_559_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	23 
    -- CP-element group 25: successors 
    -- CP-element group 25: marked-successors 
    -- CP-element group 25: 	23 
    -- CP-element group 25:  members (4) 
      -- CP-element group 25: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/ADD_u64_u64_210_sample_completed__ps
      -- CP-element group 25: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/ADD_u64_u64_210_Sample/ra
      -- CP-element group 25: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/ADD_u64_u64_210_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/ADD_u64_u64_210_sample_completed_
      -- 
    ra_618_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_210_inst_ack_0, ack => timerDaemon_CP_559_elements(25)); -- 
    -- CP-element group 26:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: marked-successors 
    -- CP-element group 26: 	24 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/ADD_u64_u64_210_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/ADD_u64_u64_210_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/ADD_u64_u64_210_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/ADD_u64_u64_210_update_completed__ps
      -- 
    ca_623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_210_inst_ack_1, ack => timerDaemon_CP_559_elements(26)); -- 
    -- CP-element group 27:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/type_cast_212_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/type_cast_212_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/type_cast_212_sample_completed__ps
      -- CP-element group 27: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/type_cast_212_sample_start__ps
      -- 
    -- Element group timerDaemon_CP_559_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (2) 
      -- CP-element group 28: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/type_cast_212_update_start_
      -- CP-element group 28: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/type_cast_212_update_start__ps
      -- 
    -- Element group timerDaemon_CP_559_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	30 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/type_cast_212_update_completed__ps
      -- 
    timerDaemon_CP_559_elements(29) <= timerDaemon_CP_559_elements(30);
    -- CP-element group 30:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	29 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/type_cast_212_update_completed_
      -- 
    -- Element group timerDaemon_CP_559_elements(30) is a control-delay.
    cp_element_30_delay: control_delay_element  generic map(name => " 30_delay", delay_value => 1)  port map(req => timerDaemon_CP_559_elements(28), ack => timerDaemon_CP_559_elements(30), clk => clk, reset =>reset);
    -- CP-element group 31:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	9 
    -- CP-element group 31: 	15 
    -- CP-element group 31: marked-predecessors 
    -- CP-element group 31: 	33 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (9) 
      -- CP-element group 31: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/STORE_count_214_Sample/word_access_start/word_0/rr
      -- CP-element group 31: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/STORE_count_214_Sample/word_access_start/word_0/$entry
      -- CP-element group 31: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/STORE_count_214_Sample/word_access_start/$entry
      -- CP-element group 31: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/STORE_count_214_Sample/STORE_count_214_Split/split_ack
      -- CP-element group 31: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/STORE_count_214_Sample/STORE_count_214_Split/split_req
      -- CP-element group 31: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/STORE_count_214_Sample/STORE_count_214_Split/$exit
      -- CP-element group 31: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/STORE_count_214_Sample/STORE_count_214_Split/$entry
      -- CP-element group 31: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/STORE_count_214_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/STORE_count_214_sample_start_
      -- 
    rr_653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_559_elements(31), ack => STORE_count_214_store_0_req_0); -- 
    timerDaemon_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 3,1 => 3,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_559_elements(9) & timerDaemon_CP_559_elements(15) & timerDaemon_CP_559_elements(33);
      gj_timerDaemon_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_559_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	34 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (5) 
      -- CP-element group 32: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/STORE_count_214_Update/word_access_complete/word_0/cr
      -- CP-element group 32: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/STORE_count_214_Update/word_access_complete/word_0/$entry
      -- CP-element group 32: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/STORE_count_214_Update/word_access_complete/$entry
      -- CP-element group 32: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/STORE_count_214_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/STORE_count_214_update_start_
      -- 
    cr_664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_559_elements(32), ack => STORE_count_214_store_0_req_1); -- 
    timerDaemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= timerDaemon_CP_559_elements(34);
      gj_timerDaemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_559_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: marked-successors 
    -- CP-element group 33: 	13 
    -- CP-element group 33: 	31 
    -- CP-element group 33:  members (5) 
      -- CP-element group 33: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/STORE_count_214_Sample/word_access_start/word_0/ra
      -- CP-element group 33: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/STORE_count_214_Sample/word_access_start/word_0/$exit
      -- CP-element group 33: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/STORE_count_214_Sample/word_access_start/$exit
      -- CP-element group 33: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/STORE_count_214_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/STORE_count_214_sample_completed_
      -- 
    ra_654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_count_214_store_0_ack_0, ack => timerDaemon_CP_559_elements(33)); -- 
    -- CP-element group 34:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34: marked-successors 
    -- CP-element group 34: 	32 
    -- CP-element group 34:  members (5) 
      -- CP-element group 34: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/STORE_count_214_Update/word_access_complete/word_0/ca
      -- CP-element group 34: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/STORE_count_214_Update/word_access_complete/word_0/$exit
      -- CP-element group 34: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/STORE_count_214_Update/word_access_complete/$exit
      -- CP-element group 34: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/STORE_count_214_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/STORE_count_214_update_completed_
      -- 
    ca_665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_count_214_store_0_ack_1, ack => timerDaemon_CP_559_elements(34)); -- 
    -- CP-element group 35:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	9 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	10 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group timerDaemon_CP_559_elements(35) is a control-delay.
    cp_element_35_delay: control_delay_element  generic map(name => " 35_delay", delay_value => 1)  port map(req => timerDaemon_CP_559_elements(9), ack => timerDaemon_CP_559_elements(35), clk => clk, reset =>reset);
    -- CP-element group 36:  join  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	14 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	6 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_203/do_while_stmt_204/do_while_stmt_204_loop_body/$exit
      -- 
    timerDaemon_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 3);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_559_elements(14) & timerDaemon_CP_559_elements(34);
      gj_timerDaemon_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_559_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	5 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (2) 
      -- CP-element group 37: 	 branch_block_stmt_203/do_while_stmt_204/loop_exit/ack
      -- CP-element group 37: 	 branch_block_stmt_203/do_while_stmt_204/loop_exit/$exit
      -- 
    ack_670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_204_branch_ack_0, ack => timerDaemon_CP_559_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	5 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (2) 
      -- CP-element group 38: 	 branch_block_stmt_203/do_while_stmt_204/loop_taken/$exit
      -- CP-element group 38: 	 branch_block_stmt_203/do_while_stmt_204/loop_taken/ack
      -- 
    ack_674_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_204_branch_ack_1, ack => timerDaemon_CP_559_elements(38)); -- 
    -- CP-element group 39:  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	3 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	1 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_203/do_while_stmt_204/$exit
      -- 
    timerDaemon_CP_559_elements(39) <= timerDaemon_CP_559_elements(3);
    timerDaemon_do_while_stmt_204_terminator_675: loop_terminator -- 
      generic map (name => " timerDaemon_do_while_stmt_204_terminator_675", max_iterations_in_flight =>3) 
      port map(loop_body_exit => timerDaemon_CP_559_elements(6),loop_continue => timerDaemon_CP_559_elements(38),loop_terminate => timerDaemon_CP_559_elements(37),loop_back => timerDaemon_CP_559_elements(4),loop_exit => timerDaemon_CP_559_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_206_phi_seq_632_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= timerDaemon_CP_559_elements(16);
      timerDaemon_CP_559_elements(21)<= src_sample_reqs(0);
      src_sample_acks(0)  <= timerDaemon_CP_559_elements(25);
      timerDaemon_CP_559_elements(22)<= src_update_reqs(0);
      src_update_acks(0)  <= timerDaemon_CP_559_elements(26);
      timerDaemon_CP_559_elements(17) <= phi_mux_reqs(0);
      triggers(1)  <= timerDaemon_CP_559_elements(18);
      timerDaemon_CP_559_elements(27)<= src_sample_reqs(1);
      src_sample_acks(1)  <= timerDaemon_CP_559_elements(27);
      timerDaemon_CP_559_elements(28)<= src_update_reqs(1);
      src_update_acks(1)  <= timerDaemon_CP_559_elements(29);
      timerDaemon_CP_559_elements(19) <= phi_mux_reqs(1);
      phi_stmt_206_phi_seq_632 : phi_sequencer_v2-- 
        generic map (place_capacity => 3, ntriggers => 2, name => "phi_stmt_206_phi_seq_632") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => timerDaemon_CP_559_elements(11), 
          phi_sample_ack => timerDaemon_CP_559_elements(14), 
          phi_update_req => timerDaemon_CP_559_elements(13), 
          phi_update_ack => timerDaemon_CP_559_elements(15), 
          phi_mux_ack => timerDaemon_CP_559_elements(20), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_584_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= timerDaemon_CP_559_elements(7);
        preds(1)  <= timerDaemon_CP_559_elements(8);
        entry_tmerge_584 : transition_merge -- 
          generic map(name => " entry_tmerge_584")
          port map (preds => preds, symbol_out => timerDaemon_CP_559_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u64_u64_210_wire : std_logic_vector(63 downto 0);
    signal STORE_count_214_data_0 : std_logic_vector(63 downto 0);
    signal STORE_count_214_word_address_0 : std_logic_vector(0 downto 0);
    signal konst_209_wire_constant : std_logic_vector(63 downto 0);
    signal konst_218_wire_constant : std_logic_vector(0 downto 0);
    signal ncount_206 : std_logic_vector(63 downto 0);
    signal type_cast_212_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    STORE_count_214_word_address_0 <= "0";
    konst_209_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_218_wire_constant <= "1";
    type_cast_212_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_206: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= ADD_u64_u64_210_wire & type_cast_212_wire_constant;
      req <= phi_stmt_206_req_0 & phi_stmt_206_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_206",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_206_ack_0,
          idata => idata,
          odata => ncount_206,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_206
    -- equivalence STORE_count_214_gather_scatter
    process(ncount_206) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ncount_206;
      ov(63 downto 0) := iv;
      STORE_count_214_data_0 <= ov(63 downto 0);
      --
    end process;
    do_while_stmt_204_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_218_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_204_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_204_branch_req_0,
          ack0 => do_while_stmt_204_branch_ack_0,
          ack1 => do_while_stmt_204_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u64_u64_210_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ncount_206;
      ADD_u64_u64_210_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_210_inst_req_0;
      ADD_u64_u64_210_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_210_inst_req_1;
      ADD_u64_u64_210_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000001",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared store operator group (0) : STORE_count_214_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 3);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_count_214_store_0_req_0;
      STORE_count_214_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_count_214_store_0_req_1;
      STORE_count_214_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_count_214_word_address_0;
      data_in <= STORE_count_214_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(0 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end timerDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity zeropad3D is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
    zeropad_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    zeropad_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    zeropad_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    zeropad_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    sendOutput_call_reqs : out  std_logic_vector(0 downto 0);
    sendOutput_call_acks : in   std_logic_vector(0 downto 0);
    sendOutput_call_data : out  std_logic_vector(31 downto 0);
    sendOutput_call_tag  :  out  std_logic_vector(0 downto 0);
    sendOutput_return_reqs : out  std_logic_vector(0 downto 0);
    sendOutput_return_acks : in   std_logic_vector(0 downto 0);
    sendOutput_return_tag :  in   std_logic_vector(0 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity zeropad3D;
architecture zeropad3D_arch of zeropad3D is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal zeropad3D_CP_676_start: Boolean;
  signal zeropad3D_CP_676_symbol: Boolean;
  -- volatile/operator module components. 
  component sendOutput is -- 
    generic (tag_length : integer); 
    port ( -- 
      size : in  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      zeropad_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal if_stmt_1331_branch_req_0 : boolean;
  signal type_cast_304_inst_req_0 : boolean;
  signal type_cast_304_inst_ack_0 : boolean;
  signal type_cast_717_inst_ack_0 : boolean;
  signal type_cast_254_inst_req_1 : boolean;
  signal W_jx_x1_761_delayed_1_0_765_inst_req_1 : boolean;
  signal phi_stmt_714_req_0 : boolean;
  signal type_cast_938_inst_req_0 : boolean;
  signal type_cast_712_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_230_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_227_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_227_inst_req_1 : boolean;
  signal type_cast_712_inst_req_1 : boolean;
  signal type_cast_266_inst_ack_0 : boolean;
  signal type_cast_653_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_230_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_227_inst_ack_0 : boolean;
  signal W_kx_x1_748_delayed_1_0_749_inst_ack_1 : boolean;
  signal type_cast_266_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_236_inst_ack_0 : boolean;
  signal ptr_deref_610_store_0_ack_1 : boolean;
  signal W_ifx_xend214_exec_guard_978_delayed_1_0_1059_inst_ack_0 : boolean;
  signal type_cast_649_inst_req_0 : boolean;
  signal type_cast_649_inst_ack_0 : boolean;
  signal type_cast_645_inst_ack_1 : boolean;
  signal phi_stmt_709_req_1 : boolean;
  signal W_lorx_xlhsx_xfalse269_exec_guard_1017_delayed_1_0_1119_inst_req_1 : boolean;
  signal type_cast_717_inst_ack_1 : boolean;
  signal type_cast_722_inst_req_0 : boolean;
  signal ptr_deref_610_store_0_req_1 : boolean;
  signal type_cast_722_inst_ack_0 : boolean;
  signal type_cast_712_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_230_inst_ack_1 : boolean;
  signal type_cast_712_inst_ack_0 : boolean;
  signal type_cast_645_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_227_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_236_inst_ack_1 : boolean;
  signal type_cast_930_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_224_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_236_inst_req_1 : boolean;
  signal type_cast_1299_inst_ack_1 : boolean;
  signal type_cast_649_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_224_inst_req_0 : boolean;
  signal type_cast_653_inst_ack_0 : boolean;
  signal W_ifx_xthen_ifx_xend214_taken_866_delayed_3_0_925_inst_ack_1 : boolean;
  signal phi_stmt_709_req_0 : boolean;
  signal type_cast_727_inst_req_1 : boolean;
  signal type_cast_1064_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_312_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_312_inst_ack_1 : boolean;
  signal phi_stmt_714_req_1 : boolean;
  signal type_cast_291_inst_req_0 : boolean;
  signal type_cast_291_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_236_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_233_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_233_inst_req_1 : boolean;
  signal type_cast_649_inst_ack_1 : boolean;
  signal type_cast_722_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_224_inst_ack_1 : boolean;
  signal type_cast_1108_inst_ack_0 : boolean;
  signal type_cast_266_inst_ack_1 : boolean;
  signal W_jx_x1_761_delayed_1_0_765_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_287_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_287_inst_ack_0 : boolean;
  signal W_lorx_xlhsx_xfalse269_exec_guard_1017_delayed_1_0_1119_inst_ack_1 : boolean;
  signal type_cast_279_inst_req_1 : boolean;
  signal type_cast_279_inst_ack_0 : boolean;
  signal type_cast_279_inst_req_0 : boolean;
  signal W_kx_x1_748_delayed_1_0_749_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_275_inst_req_0 : boolean;
  signal type_cast_241_inst_ack_1 : boolean;
  signal type_cast_241_inst_req_1 : boolean;
  signal type_cast_1347_inst_req_1 : boolean;
  signal ptr_deref_1268_load_0_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_262_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_262_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_262_inst_ack_0 : boolean;
  signal type_cast_645_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_250_inst_req_0 : boolean;
  signal type_cast_254_inst_ack_0 : boolean;
  signal type_cast_254_inst_req_0 : boolean;
  signal W_ifx_xthen_ifx_xend214_taken_882_delayed_3_0_953_inst_ack_1 : boolean;
  signal phi_stmt_709_ack_0 : boolean;
  signal type_cast_1277_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_262_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_275_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_287_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_287_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_275_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_230_inst_req_1 : boolean;
  signal type_cast_241_inst_ack_0 : boolean;
  signal type_cast_241_inst_req_0 : boolean;
  signal type_cast_722_inst_ack_1 : boolean;
  signal W_jx_x1_761_delayed_1_0_765_inst_ack_0 : boolean;
  signal type_cast_266_inst_req_1 : boolean;
  signal type_cast_291_inst_req_1 : boolean;
  signal type_cast_291_inst_ack_1 : boolean;
  signal type_cast_254_inst_ack_1 : boolean;
  signal type_cast_304_inst_req_1 : boolean;
  signal type_cast_304_inst_ack_1 : boolean;
  signal type_cast_717_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_312_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_312_inst_ack_0 : boolean;
  signal type_cast_778_inst_ack_1 : boolean;
  signal type_cast_653_inst_req_0 : boolean;
  signal type_cast_1064_inst_req_0 : boolean;
  signal type_cast_279_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_300_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_300_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_250_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_233_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_300_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_300_inst_ack_0 : boolean;
  signal call_stmt_635_call_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_250_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_233_inst_req_0 : boolean;
  signal type_cast_727_inst_ack_1 : boolean;
  signal call_stmt_635_call_req_1 : boolean;
  signal type_cast_645_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_275_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_250_inst_ack_0 : boolean;
  signal type_cast_653_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_224_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_315_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_315_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_315_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_315_inst_ack_1 : boolean;
  signal type_cast_934_inst_ack_1 : boolean;
  signal type_cast_717_inst_req_0 : boolean;
  signal phi_stmt_719_ack_0 : boolean;
  signal type_cast_319_inst_req_0 : boolean;
  signal type_cast_319_inst_ack_0 : boolean;
  signal type_cast_319_inst_req_1 : boolean;
  signal type_cast_319_inst_ack_1 : boolean;
  signal type_cast_778_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_328_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_328_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_328_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_328_inst_ack_1 : boolean;
  signal W_ifx_xthen_ifx_xend214_taken_866_delayed_3_0_925_inst_req_0 : boolean;
  signal W_add230_1128_delayed_2_0_1270_inst_ack_1 : boolean;
  signal type_cast_332_inst_req_0 : boolean;
  signal type_cast_332_inst_ack_0 : boolean;
  signal type_cast_332_inst_req_1 : boolean;
  signal type_cast_332_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_340_inst_req_0 : boolean;
  signal type_cast_1038_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_340_inst_ack_0 : boolean;
  signal call_stmt_635_call_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_340_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_340_inst_ack_1 : boolean;
  signal W_ifx_xend214_exec_guard_978_delayed_1_0_1059_inst_req_0 : boolean;
  signal type_cast_344_inst_req_0 : boolean;
  signal type_cast_344_inst_ack_0 : boolean;
  signal type_cast_344_inst_req_1 : boolean;
  signal type_cast_344_inst_ack_1 : boolean;
  signal type_cast_727_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_353_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_353_inst_ack_0 : boolean;
  signal call_stmt_635_call_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_353_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_353_inst_ack_1 : boolean;
  signal type_cast_934_inst_req_0 : boolean;
  signal type_cast_357_inst_req_0 : boolean;
  signal type_cast_357_inst_ack_0 : boolean;
  signal type_cast_357_inst_req_1 : boolean;
  signal type_cast_357_inst_ack_1 : boolean;
  signal type_cast_727_inst_req_0 : boolean;
  signal type_cast_778_inst_ack_0 : boolean;
  signal W_ifx_xthen_ifx_xend214_taken_866_delayed_3_0_925_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_365_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_365_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_365_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_365_inst_ack_1 : boolean;
  signal W_lorx_xlhsx_xfalse269_exec_guard_1039_delayed_1_0_1152_inst_ack_1 : boolean;
  signal array_obj_ref_1305_index_offset_ack_0 : boolean;
  signal type_cast_1038_inst_req_1 : boolean;
  signal type_cast_938_inst_req_1 : boolean;
  signal type_cast_1038_inst_ack_1 : boolean;
  signal type_cast_369_inst_req_0 : boolean;
  signal type_cast_369_inst_ack_0 : boolean;
  signal type_cast_369_inst_req_1 : boolean;
  signal type_cast_369_inst_ack_1 : boolean;
  signal type_cast_778_inst_req_0 : boolean;
  signal W_ifx_xend214_exec_guard_971_delayed_1_0_1049_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_378_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_378_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_378_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_378_inst_ack_1 : boolean;
  signal ptr_deref_610_store_0_ack_0 : boolean;
  signal type_cast_382_inst_req_0 : boolean;
  signal type_cast_382_inst_ack_0 : boolean;
  signal type_cast_382_inst_req_1 : boolean;
  signal type_cast_382_inst_ack_1 : boolean;
  signal type_cast_938_inst_ack_1 : boolean;
  signal type_cast_391_inst_req_0 : boolean;
  signal type_cast_391_inst_ack_0 : boolean;
  signal W_ifx_xend214_exec_guard_993_delayed_1_0_1082_inst_req_1 : boolean;
  signal phi_stmt_719_req_1 : boolean;
  signal type_cast_391_inst_req_1 : boolean;
  signal type_cast_391_inst_ack_1 : boolean;
  signal type_cast_938_inst_ack_0 : boolean;
  signal type_cast_395_inst_req_0 : boolean;
  signal type_cast_395_inst_ack_0 : boolean;
  signal type_cast_395_inst_req_1 : boolean;
  signal type_cast_395_inst_ack_1 : boolean;
  signal type_cast_399_inst_req_0 : boolean;
  signal type_cast_399_inst_ack_0 : boolean;
  signal W_ifx_xend214_exec_guard_993_delayed_1_0_1082_inst_ack_1 : boolean;
  signal W_add230_1128_delayed_2_0_1270_inst_req_0 : boolean;
  signal type_cast_399_inst_req_1 : boolean;
  signal type_cast_399_inst_ack_1 : boolean;
  signal W_ifx_xthen_ifx_xend214_taken_882_delayed_3_0_953_inst_req_1 : boolean;
  signal type_cast_934_inst_req_1 : boolean;
  signal W_kx_x1_748_delayed_1_0_749_inst_ack_0 : boolean;
  signal W_ifx_xthen_ifx_xend214_taken_866_delayed_3_0_925_inst_ack_0 : boolean;
  signal W_ifx_xend214_exec_guard_978_delayed_1_0_1059_inst_req_1 : boolean;
  signal ptr_deref_610_store_0_req_0 : boolean;
  signal W_ifx_xend214_exec_guard_993_delayed_1_0_1082_inst_req_0 : boolean;
  signal if_stmt_433_branch_req_0 : boolean;
  signal do_while_stmt_707_branch_req_0 : boolean;
  signal if_stmt_433_branch_ack_1 : boolean;
  signal if_stmt_433_branch_ack_0 : boolean;
  signal W_ifx_xend214_exec_guard_978_delayed_1_0_1059_inst_ack_1 : boolean;
  signal phi_stmt_714_ack_0 : boolean;
  signal array_obj_ref_1305_index_offset_req_0 : boolean;
  signal type_cast_731_inst_ack_1 : boolean;
  signal array_obj_ref_473_index_offset_req_0 : boolean;
  signal array_obj_ref_473_index_offset_ack_0 : boolean;
  signal type_cast_731_inst_req_1 : boolean;
  signal array_obj_ref_473_index_offset_req_1 : boolean;
  signal array_obj_ref_473_index_offset_ack_1 : boolean;
  signal W_jx_x1_761_delayed_1_0_765_inst_ack_1 : boolean;
  signal W_kx_x1_748_delayed_1_0_749_inst_req_0 : boolean;
  signal type_cast_1038_inst_ack_0 : boolean;
  signal addr_of_474_final_reg_req_0 : boolean;
  signal addr_of_474_final_reg_ack_0 : boolean;
  signal W_ifx_xend214_exec_guard_993_delayed_1_0_1082_inst_ack_0 : boolean;
  signal addr_of_474_final_reg_req_1 : boolean;
  signal addr_of_474_final_reg_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_477_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_477_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_477_inst_req_1 : boolean;
  signal W_arrayidx303_1156_delayed_5_0_1311_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_477_inst_ack_1 : boolean;
  signal type_cast_677_inst_ack_1 : boolean;
  signal type_cast_677_inst_req_1 : boolean;
  signal phi_stmt_719_req_0 : boolean;
  signal type_cast_481_inst_req_0 : boolean;
  signal type_cast_481_inst_ack_0 : boolean;
  signal type_cast_930_inst_req_1 : boolean;
  signal type_cast_481_inst_req_1 : boolean;
  signal type_cast_481_inst_ack_1 : boolean;
  signal if_stmt_624_branch_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_490_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_490_inst_ack_0 : boolean;
  signal type_cast_731_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_490_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_490_inst_ack_1 : boolean;
  signal type_cast_677_inst_ack_0 : boolean;
  signal type_cast_1299_inst_req_1 : boolean;
  signal type_cast_677_inst_req_0 : boolean;
  signal type_cast_494_inst_req_0 : boolean;
  signal type_cast_494_inst_ack_0 : boolean;
  signal type_cast_494_inst_req_1 : boolean;
  signal type_cast_494_inst_ack_1 : boolean;
  signal if_stmt_624_branch_ack_1 : boolean;
  signal type_cast_731_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_508_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_508_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_508_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_508_inst_ack_1 : boolean;
  signal type_cast_668_inst_ack_1 : boolean;
  signal type_cast_668_inst_req_1 : boolean;
  signal type_cast_668_inst_ack_0 : boolean;
  signal type_cast_668_inst_req_0 : boolean;
  signal type_cast_512_inst_req_0 : boolean;
  signal type_cast_512_inst_ack_0 : boolean;
  signal type_cast_512_inst_req_1 : boolean;
  signal type_cast_512_inst_ack_1 : boolean;
  signal if_stmt_624_branch_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_526_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_526_inst_ack_0 : boolean;
  signal W_arrayidx303_1156_delayed_5_0_1311_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_526_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_526_inst_ack_1 : boolean;
  signal type_cast_530_inst_req_0 : boolean;
  signal type_cast_530_inst_ack_0 : boolean;
  signal type_cast_530_inst_req_1 : boolean;
  signal type_cast_530_inst_ack_1 : boolean;
  signal W_ifx_xthen_ifx_xend214_taken_882_delayed_3_0_953_inst_req_0 : boolean;
  signal type_cast_1064_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_544_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_544_inst_ack_0 : boolean;
  signal type_cast_930_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_544_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_544_inst_ack_1 : boolean;
  signal do_while_stmt_707_branch_ack_1 : boolean;
  signal type_cast_548_inst_req_0 : boolean;
  signal type_cast_1064_inst_ack_1 : boolean;
  signal type_cast_548_inst_ack_0 : boolean;
  signal type_cast_548_inst_req_1 : boolean;
  signal type_cast_548_inst_ack_1 : boolean;
  signal W_ifx_xthen_ifx_xend214_taken_882_delayed_3_0_953_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_562_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_562_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_562_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_562_inst_ack_1 : boolean;
  signal type_cast_930_inst_ack_0 : boolean;
  signal type_cast_566_inst_req_0 : boolean;
  signal type_cast_566_inst_ack_0 : boolean;
  signal type_cast_1108_inst_req_0 : boolean;
  signal type_cast_566_inst_req_1 : boolean;
  signal type_cast_566_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_580_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_580_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_580_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_580_inst_ack_1 : boolean;
  signal type_cast_584_inst_req_0 : boolean;
  signal type_cast_584_inst_ack_0 : boolean;
  signal type_cast_584_inst_req_1 : boolean;
  signal type_cast_584_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_598_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_598_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_598_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_598_inst_ack_1 : boolean;
  signal type_cast_602_inst_req_0 : boolean;
  signal type_cast_602_inst_ack_0 : boolean;
  signal type_cast_602_inst_req_1 : boolean;
  signal type_cast_602_inst_ack_1 : boolean;
  signal W_lorx_xlhsx_xfalse269_exec_guard_1039_delayed_1_0_1152_inst_ack_0 : boolean;
  signal W_ifx_xend214_exec_guard_971_delayed_1_0_1049_inst_req_1 : boolean;
  signal W_lorx_xlhsx_xfalse269_exec_guard_1017_delayed_1_0_1119_inst_ack_0 : boolean;
  signal W_ifx_xelse_exec_guard_771_delayed_1_0_780_inst_req_0 : boolean;
  signal W_ifx_xelse_exec_guard_771_delayed_1_0_780_inst_ack_0 : boolean;
  signal type_cast_1299_inst_req_0 : boolean;
  signal W_ifx_xelse_exec_guard_771_delayed_1_0_780_inst_req_1 : boolean;
  signal W_ifx_xelse_exec_guard_771_delayed_1_0_780_inst_ack_1 : boolean;
  signal W_lorx_xlhsx_xfalse269_exec_guard_1017_delayed_1_0_1119_inst_req_0 : boolean;
  signal W_ifx_xelse_exec_guard_777_delayed_1_0_789_inst_req_0 : boolean;
  signal W_ifx_xend214_exec_guard_998_delayed_1_0_1090_inst_ack_1 : boolean;
  signal W_ifx_xelse_exec_guard_777_delayed_1_0_789_inst_ack_0 : boolean;
  signal W_ifx_xelse_exec_guard_777_delayed_1_0_789_inst_req_1 : boolean;
  signal W_ifx_xelse_exec_guard_777_delayed_1_0_789_inst_ack_1 : boolean;
  signal ptr_deref_1316_store_0_req_1 : boolean;
  signal W_lorx_xlhsx_xfalse269_exec_guard_1039_delayed_1_0_1152_inst_req_0 : boolean;
  signal W_ifx_xend214_exec_guard_998_delayed_1_0_1090_inst_req_1 : boolean;
  signal type_cast_795_inst_req_0 : boolean;
  signal type_cast_795_inst_ack_0 : boolean;
  signal W_ifx_xend214_exec_guard_986_delayed_1_0_1073_inst_ack_1 : boolean;
  signal type_cast_795_inst_req_1 : boolean;
  signal type_cast_795_inst_ack_1 : boolean;
  signal type_cast_1366_inst_req_0 : boolean;
  signal W_ifx_xend214_exec_guard_971_delayed_1_0_1049_inst_ack_0 : boolean;
  signal W_ifx_xelse_exec_guard_782_delayed_2_0_797_inst_req_0 : boolean;
  signal W_ifx_xelse_exec_guard_782_delayed_2_0_797_inst_ack_0 : boolean;
  signal W_ifx_xelse_exec_guard_782_delayed_2_0_797_inst_req_1 : boolean;
  signal W_ifx_xelse_exec_guard_782_delayed_2_0_797_inst_ack_1 : boolean;
  signal type_cast_1356_inst_req_0 : boolean;
  signal W_ifx_xend214_exec_guard_971_delayed_1_0_1049_inst_req_0 : boolean;
  signal W_i138x_x2_785_delayed_3_0_800_inst_req_0 : boolean;
  signal W_ifx_xend214_exec_guard_998_delayed_1_0_1090_inst_ack_0 : boolean;
  signal W_i138x_x2_785_delayed_3_0_800_inst_ack_0 : boolean;
  signal type_cast_1299_inst_ack_0 : boolean;
  signal W_i138x_x2_785_delayed_3_0_800_inst_req_1 : boolean;
  signal W_i138x_x2_785_delayed_3_0_800_inst_ack_1 : boolean;
  signal type_cast_1347_inst_req_0 : boolean;
  signal type_cast_1277_inst_ack_1 : boolean;
  signal ptr_deref_1268_load_0_req_0 : boolean;
  signal W_ifx_xelse_exec_guard_788_delayed_1_0_809_inst_req_0 : boolean;
  signal W_ifx_xend214_exec_guard_998_delayed_1_0_1090_inst_req_0 : boolean;
  signal W_ifx_xelse_exec_guard_788_delayed_1_0_809_inst_ack_0 : boolean;
  signal W_add230_1128_delayed_2_0_1270_inst_ack_0 : boolean;
  signal W_ifx_xelse_exec_guard_788_delayed_1_0_809_inst_req_1 : boolean;
  signal W_ifx_xelse_exec_guard_788_delayed_1_0_809_inst_ack_1 : boolean;
  signal W_lorx_xlhsx_xfalse269_exec_guard_1044_delayed_1_0_1160_inst_ack_1 : boolean;
  signal W_lorx_xlhsx_xfalse269_exec_guard_1039_delayed_1_0_1152_inst_req_1 : boolean;
  signal W_ifx_xend214_ifx_xthen286_taken_1050_delayed_1_0_1169_inst_ack_1 : boolean;
  signal W_inc187_793_delayed_1_0_812_inst_req_0 : boolean;
  signal W_inc187_793_delayed_1_0_812_inst_ack_0 : boolean;
  signal W_inc187_793_delayed_1_0_812_inst_req_1 : boolean;
  signal W_inc187_793_delayed_1_0_812_inst_ack_1 : boolean;
  signal type_cast_1356_inst_ack_0 : boolean;
  signal W_lorx_xlhsx_xfalse269_exec_guard_1044_delayed_1_0_1160_inst_req_1 : boolean;
  signal type_cast_1347_inst_ack_0 : boolean;
  signal type_cast_1386_inst_req_1 : boolean;
  signal type_cast_1108_inst_ack_1 : boolean;
  signal W_ifx_xelse_exec_guard_796_delayed_2_0_823_inst_req_0 : boolean;
  signal W_arrayidx303_1156_delayed_5_0_1311_inst_req_1 : boolean;
  signal W_ifx_xelse_exec_guard_796_delayed_2_0_823_inst_ack_0 : boolean;
  signal W_ifx_xelse_exec_guard_796_delayed_2_0_823_inst_req_1 : boolean;
  signal W_ifx_xelse_exec_guard_796_delayed_2_0_823_inst_ack_1 : boolean;
  signal do_while_stmt_707_branch_ack_0 : boolean;
  signal W_ifx_xend214_ifx_xthen286_taken_1050_delayed_1_0_1169_inst_req_1 : boolean;
  signal W_ifx_xelse292_exec_guard_1155_delayed_14_0_1308_inst_ack_1 : boolean;
  signal W_add230_1128_delayed_2_0_1270_inst_req_1 : boolean;
  signal W_jx_x0_1008_delayed_1_0_1102_inst_ack_1 : boolean;
  signal if_stmt_1331_branch_ack_1 : boolean;
  signal type_cast_1108_inst_req_1 : boolean;
  signal W_jx_x0_1008_delayed_1_0_1102_inst_req_1 : boolean;
  signal type_cast_829_inst_req_0 : boolean;
  signal type_cast_829_inst_ack_0 : boolean;
  signal W_ifx_xend214_exec_guard_986_delayed_1_0_1073_inst_req_1 : boolean;
  signal type_cast_829_inst_req_1 : boolean;
  signal type_cast_829_inst_ack_1 : boolean;
  signal W_ifx_xelse_exec_guard_801_delayed_3_0_831_inst_req_0 : boolean;
  signal W_ifx_xelse_exec_guard_801_delayed_3_0_831_inst_ack_0 : boolean;
  signal W_ifx_xelse_exec_guard_801_delayed_3_0_831_inst_req_1 : boolean;
  signal W_ifx_xelse_exec_guard_801_delayed_3_0_831_inst_ack_1 : boolean;
  signal W_lorx_xlhsx_xfalse269_exec_guard_1044_delayed_1_0_1160_inst_ack_0 : boolean;
  signal W_ifx_xelse_exec_guard_808_delayed_3_0_840_inst_req_0 : boolean;
  signal W_ifx_xelse_exec_guard_808_delayed_3_0_840_inst_ack_0 : boolean;
  signal W_ifx_xelse_exec_guard_808_delayed_3_0_840_inst_req_1 : boolean;
  signal W_arrayidx303_1156_delayed_5_0_1311_inst_ack_1 : boolean;
  signal W_ifx_xelse_exec_guard_808_delayed_3_0_840_inst_ack_1 : boolean;
  signal W_lorx_xlhsx_xfalse269_exec_guard_1044_delayed_1_0_1160_inst_req_0 : boolean;
  signal W_jx_x0_1008_delayed_1_0_1102_inst_ack_0 : boolean;
  signal W_ifx_xelse_exec_guard_813_delayed_3_0_848_inst_req_0 : boolean;
  signal W_ifx_xelse_exec_guard_813_delayed_3_0_848_inst_ack_0 : boolean;
  signal W_ifx_xelse_exec_guard_813_delayed_3_0_848_inst_req_1 : boolean;
  signal W_ifx_xelse_exec_guard_813_delayed_3_0_848_inst_ack_1 : boolean;
  signal W_lorx_xlhsx_xfalse269_exec_guard_1032_delayed_1_0_1143_inst_ack_1 : boolean;
  signal W_lorx_xlhsx_xfalse269_exec_guard_1024_delayed_1_0_1129_inst_ack_1 : boolean;
  signal W_lorx_xlhsx_xfalse269_exec_guard_1024_delayed_1_0_1129_inst_req_1 : boolean;
  signal type_cast_1134_inst_ack_0 : boolean;
  signal W_ifx_xend214_ifx_xthen286_taken_1050_delayed_1_0_1169_inst_ack_0 : boolean;
  signal W_jx_x0_1008_delayed_1_0_1102_inst_req_0 : boolean;
  signal W_ifx_xend214_exec_guard_965_delayed_1_0_1040_inst_ack_1 : boolean;
  signal W_ifx_xthen_ifx_xend214_taken_826_delayed_3_0_863_inst_req_0 : boolean;
  signal W_ifx_xthen_ifx_xend214_taken_826_delayed_3_0_863_inst_ack_0 : boolean;
  signal W_ifx_xthen_ifx_xend214_taken_826_delayed_3_0_863_inst_req_1 : boolean;
  signal W_ifx_xthen_ifx_xend214_taken_826_delayed_3_0_863_inst_ack_1 : boolean;
  signal W_lorx_xlhsx_xfalse269_exec_guard_1032_delayed_1_0_1143_inst_req_1 : boolean;
  signal type_cast_1134_inst_req_0 : boolean;
  signal W_ifx_xend214_ifx_xthen286_taken_1050_delayed_1_0_1169_inst_req_0 : boolean;
  signal type_cast_1386_inst_req_0 : boolean;
  signal W_ifx_xend214_exec_guard_965_delayed_1_0_1040_inst_req_1 : boolean;
  signal W_ifx_xthen_ifx_xend214_taken_832_delayed_3_0_873_inst_req_0 : boolean;
  signal W_ifx_xthen_ifx_xend214_taken_832_delayed_3_0_873_inst_ack_0 : boolean;
  signal W_ifx_xthen_ifx_xend214_taken_832_delayed_3_0_873_inst_req_1 : boolean;
  signal W_ifx_xthen_ifx_xend214_taken_832_delayed_3_0_873_inst_ack_1 : boolean;
  signal W_lorx_xlhsx_xfalse269_exec_guard_1024_delayed_1_0_1129_inst_ack_0 : boolean;
  signal type_cast_878_inst_req_0 : boolean;
  signal type_cast_878_inst_ack_0 : boolean;
  signal type_cast_878_inst_req_1 : boolean;
  signal type_cast_878_inst_ack_1 : boolean;
  signal ptr_deref_1316_store_0_ack_1 : boolean;
  signal W_lorx_xlhsx_xfalse269_exec_guard_1024_delayed_1_0_1129_inst_req_0 : boolean;
  signal W_ifx_xelse292_exec_guard_1142_delayed_1_0_1292_inst_req_1 : boolean;
  signal type_cast_1386_inst_ack_0 : boolean;
  signal type_cast_1396_inst_ack_0 : boolean;
  signal W_ifx_xelse292_exec_guard_1142_delayed_1_0_1292_inst_ack_0 : boolean;
  signal W_ifx_xend214_exec_guard_965_delayed_1_0_1040_inst_ack_0 : boolean;
  signal W_lorx_xlhsx_xfalse269_exec_guard_1011_delayed_1_0_1110_inst_ack_1 : boolean;
  signal W_ifx_xthen_ifx_xend214_taken_850_delayed_3_0_897_inst_req_0 : boolean;
  signal W_ifx_xthen_ifx_xend214_taken_850_delayed_3_0_897_inst_ack_0 : boolean;
  signal W_ifx_xthen_ifx_xend214_taken_850_delayed_3_0_897_inst_req_1 : boolean;
  signal W_ifx_xthen_ifx_xend214_taken_850_delayed_3_0_897_inst_ack_1 : boolean;
  signal W_lorx_xlhsx_xfalse269_exec_guard_1032_delayed_1_0_1143_inst_ack_0 : boolean;
  signal type_cast_1134_inst_ack_1 : boolean;
  signal W_lorx_xlhsx_xfalse269_exec_guard_1032_delayed_1_0_1143_inst_req_0 : boolean;
  signal W_ifx_xend214_exec_guard_965_delayed_1_0_1040_inst_req_0 : boolean;
  signal W_lorx_xlhsx_xfalse269_exec_guard_1011_delayed_1_0_1110_inst_req_1 : boolean;
  signal type_cast_902_inst_req_0 : boolean;
  signal type_cast_902_inst_ack_0 : boolean;
  signal type_cast_902_inst_req_1 : boolean;
  signal type_cast_902_inst_ack_1 : boolean;
  signal if_stmt_1331_branch_ack_0 : boolean;
  signal type_cast_906_inst_req_0 : boolean;
  signal type_cast_906_inst_ack_0 : boolean;
  signal W_lorx_xlhsx_xfalse269_exec_guard_1011_delayed_1_0_1110_inst_ack_0 : boolean;
  signal type_cast_906_inst_req_1 : boolean;
  signal type_cast_906_inst_ack_1 : boolean;
  signal type_cast_1134_inst_req_1 : boolean;
  signal W_ifx_xelse292_exec_guard_1155_delayed_14_0_1308_inst_req_1 : boolean;
  signal W_ifx_xend214_exec_guard_986_delayed_1_0_1073_inst_ack_0 : boolean;
  signal W_lorx_xlhsx_xfalse269_exec_guard_1011_delayed_1_0_1110_inst_req_0 : boolean;
  signal type_cast_910_inst_req_0 : boolean;
  signal type_cast_910_inst_ack_0 : boolean;
  signal W_ifx_xend214_exec_guard_986_delayed_1_0_1073_inst_req_0 : boolean;
  signal type_cast_910_inst_req_1 : boolean;
  signal type_cast_910_inst_ack_1 : boolean;
  signal type_cast_1396_inst_req_1 : boolean;
  signal type_cast_1396_inst_ack_1 : boolean;
  signal type_cast_1366_inst_ack_0 : boolean;
  signal type_cast_1347_inst_ack_1 : boolean;
  signal W_ifx_xelse292_exec_guard_1142_delayed_1_0_1292_inst_ack_1 : boolean;
  signal type_cast_934_inst_ack_0 : boolean;
  signal W_add230_1056_delayed_2_0_1177_inst_req_0 : boolean;
  signal W_add230_1056_delayed_2_0_1177_inst_ack_0 : boolean;
  signal W_add230_1056_delayed_2_0_1177_inst_req_1 : boolean;
  signal W_add230_1056_delayed_2_0_1177_inst_ack_1 : boolean;
  signal type_cast_1396_inst_req_0 : boolean;
  signal type_cast_1366_inst_ack_1 : boolean;
  signal ptr_deref_1316_store_0_ack_0 : boolean;
  signal W_ifx_xelse292_exec_guard_1155_delayed_14_0_1308_inst_ack_0 : boolean;
  signal call_stmt_1343_call_ack_1 : boolean;
  signal type_cast_1184_inst_req_0 : boolean;
  signal W_ifx_xelse292_exec_guard_1155_delayed_14_0_1308_inst_req_0 : boolean;
  signal type_cast_1184_inst_ack_0 : boolean;
  signal call_stmt_1343_call_req_1 : boolean;
  signal type_cast_1184_inst_req_1 : boolean;
  signal type_cast_1184_inst_ack_1 : boolean;
  signal ptr_deref_1316_store_0_req_0 : boolean;
  signal W_ifx_xelse292_exec_guard_1142_delayed_1_0_1292_inst_req_0 : boolean;
  signal W_ifx_xthen286_exec_guard_1060_delayed_1_0_1186_inst_req_0 : boolean;
  signal W_ifx_xthen286_exec_guard_1060_delayed_1_0_1186_inst_ack_0 : boolean;
  signal W_ifx_xthen286_exec_guard_1060_delayed_1_0_1186_inst_req_1 : boolean;
  signal W_ifx_xthen286_exec_guard_1060_delayed_1_0_1186_inst_ack_1 : boolean;
  signal type_cast_1376_inst_ack_1 : boolean;
  signal type_cast_1366_inst_req_1 : boolean;
  signal type_cast_1376_inst_req_1 : boolean;
  signal type_cast_1376_inst_req_0 : boolean;
  signal W_ifx_xthen286_exec_guard_1070_delayed_1_0_1199_inst_req_0 : boolean;
  signal W_ifx_xthen286_exec_guard_1070_delayed_1_0_1199_inst_ack_0 : boolean;
  signal W_ifx_xthen286_exec_guard_1070_delayed_1_0_1199_inst_req_1 : boolean;
  signal W_ifx_xthen286_exec_guard_1070_delayed_1_0_1199_inst_ack_1 : boolean;
  signal call_stmt_1343_call_ack_0 : boolean;
  signal call_stmt_1343_call_req_0 : boolean;
  signal type_cast_1206_inst_req_0 : boolean;
  signal addr_of_1306_final_reg_ack_1 : boolean;
  signal type_cast_1206_inst_ack_0 : boolean;
  signal type_cast_1206_inst_req_1 : boolean;
  signal addr_of_1306_final_reg_req_1 : boolean;
  signal type_cast_1206_inst_ack_1 : boolean;
  signal W_ifx_xelse292_exec_guard_1132_delayed_1_0_1279_inst_ack_1 : boolean;
  signal array_obj_ref_1212_index_offset_req_0 : boolean;
  signal array_obj_ref_1212_index_offset_ack_0 : boolean;
  signal array_obj_ref_1212_index_offset_req_1 : boolean;
  signal array_obj_ref_1212_index_offset_ack_1 : boolean;
  signal type_cast_1339_inst_ack_1 : boolean;
  signal addr_of_1306_final_reg_ack_0 : boolean;
  signal addr_of_1306_final_reg_req_0 : boolean;
  signal addr_of_1213_final_reg_req_0 : boolean;
  signal addr_of_1213_final_reg_ack_0 : boolean;
  signal addr_of_1213_final_reg_req_1 : boolean;
  signal addr_of_1213_final_reg_ack_1 : boolean;
  signal W_ifx_xelse292_exec_guard_1132_delayed_1_0_1279_inst_req_1 : boolean;
  signal type_cast_1277_inst_ack_0 : boolean;
  signal type_cast_1277_inst_req_0 : boolean;
  signal ptr_deref_1217_store_0_req_0 : boolean;
  signal W_ifx_xelse292_exec_guard_1132_delayed_1_0_1279_inst_ack_0 : boolean;
  signal ptr_deref_1217_store_0_ack_0 : boolean;
  signal ptr_deref_1217_store_0_req_1 : boolean;
  signal W_ifx_xelse292_exec_guard_1132_delayed_1_0_1279_inst_req_0 : boolean;
  signal ptr_deref_1217_store_0_ack_1 : boolean;
  signal type_cast_1386_inst_ack_1 : boolean;
  signal type_cast_1339_inst_req_1 : boolean;
  signal W_add252_1094_delayed_2_0_1224_inst_req_0 : boolean;
  signal array_obj_ref_1305_index_offset_ack_1 : boolean;
  signal W_add252_1094_delayed_2_0_1224_inst_ack_0 : boolean;
  signal W_add252_1094_delayed_2_0_1224_inst_req_1 : boolean;
  signal array_obj_ref_1305_index_offset_req_1 : boolean;
  signal W_add252_1094_delayed_2_0_1224_inst_ack_1 : boolean;
  signal type_cast_1376_inst_ack_0 : boolean;
  signal ptr_deref_1268_load_0_ack_1 : boolean;
  signal ptr_deref_1268_load_0_req_1 : boolean;
  signal type_cast_1356_inst_ack_1 : boolean;
  signal type_cast_1356_inst_req_1 : boolean;
  signal type_cast_1339_inst_ack_0 : boolean;
  signal type_cast_1339_inst_req_0 : boolean;
  signal type_cast_1231_inst_req_0 : boolean;
  signal type_cast_1231_inst_ack_0 : boolean;
  signal type_cast_1231_inst_req_1 : boolean;
  signal type_cast_1231_inst_ack_1 : boolean;
  signal W_ifx_xelse292_exec_guard_1098_delayed_1_0_1233_inst_req_0 : boolean;
  signal W_ifx_xelse292_exec_guard_1098_delayed_1_0_1233_inst_ack_0 : boolean;
  signal W_ifx_xelse292_exec_guard_1098_delayed_1_0_1233_inst_req_1 : boolean;
  signal W_ifx_xelse292_exec_guard_1098_delayed_1_0_1233_inst_ack_1 : boolean;
  signal W_ifx_xelse292_exec_guard_1108_delayed_1_0_1246_inst_req_0 : boolean;
  signal W_ifx_xelse292_exec_guard_1108_delayed_1_0_1246_inst_ack_0 : boolean;
  signal W_ifx_xelse292_exec_guard_1108_delayed_1_0_1246_inst_req_1 : boolean;
  signal W_ifx_xelse292_exec_guard_1108_delayed_1_0_1246_inst_ack_1 : boolean;
  signal type_cast_1253_inst_req_0 : boolean;
  signal type_cast_1253_inst_ack_0 : boolean;
  signal type_cast_1253_inst_req_1 : boolean;
  signal type_cast_1253_inst_ack_1 : boolean;
  signal array_obj_ref_1259_index_offset_req_0 : boolean;
  signal array_obj_ref_1259_index_offset_ack_0 : boolean;
  signal array_obj_ref_1259_index_offset_req_1 : boolean;
  signal array_obj_ref_1259_index_offset_ack_1 : boolean;
  signal addr_of_1260_final_reg_req_0 : boolean;
  signal addr_of_1260_final_reg_ack_0 : boolean;
  signal addr_of_1260_final_reg_req_1 : boolean;
  signal addr_of_1260_final_reg_ack_1 : boolean;
  signal W_ifx_xelse292_exec_guard_1121_delayed_8_0_1262_inst_req_0 : boolean;
  signal W_ifx_xelse292_exec_guard_1121_delayed_8_0_1262_inst_ack_0 : boolean;
  signal W_ifx_xelse292_exec_guard_1121_delayed_8_0_1262_inst_req_1 : boolean;
  signal W_ifx_xelse292_exec_guard_1121_delayed_8_0_1262_inst_ack_1 : boolean;
  signal type_cast_1406_inst_req_0 : boolean;
  signal type_cast_1406_inst_ack_0 : boolean;
  signal type_cast_1406_inst_req_1 : boolean;
  signal type_cast_1406_inst_ack_1 : boolean;
  signal type_cast_1416_inst_req_0 : boolean;
  signal type_cast_1416_inst_ack_0 : boolean;
  signal type_cast_1416_inst_req_1 : boolean;
  signal type_cast_1416_inst_ack_1 : boolean;
  signal type_cast_1426_inst_req_0 : boolean;
  signal type_cast_1426_inst_ack_0 : boolean;
  signal type_cast_1426_inst_req_1 : boolean;
  signal type_cast_1426_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_1428_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_1428_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_1428_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_1428_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_1431_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_1431_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_1431_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_1431_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_1434_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_1434_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_1434_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_1434_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_1437_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_1437_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_1437_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_1437_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_1440_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_1440_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_1440_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_1440_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_1443_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_1443_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_1443_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_1443_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_1446_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_1446_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_1446_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_1446_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_1449_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_1449_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_1449_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_1449_inst_ack_1 : boolean;
  signal type_cast_1455_inst_req_0 : boolean;
  signal type_cast_1455_inst_ack_0 : boolean;
  signal type_cast_1455_inst_req_1 : boolean;
  signal type_cast_1455_inst_ack_1 : boolean;
  signal type_cast_1459_inst_req_0 : boolean;
  signal type_cast_1459_inst_ack_0 : boolean;
  signal type_cast_1459_inst_req_1 : boolean;
  signal type_cast_1459_inst_ack_1 : boolean;
  signal call_stmt_1472_call_req_0 : boolean;
  signal call_stmt_1472_call_ack_0 : boolean;
  signal call_stmt_1472_call_req_1 : boolean;
  signal call_stmt_1472_call_ack_1 : boolean;
  signal phi_stmt_461_req_0 : boolean;
  signal type_cast_467_inst_req_0 : boolean;
  signal type_cast_467_inst_ack_0 : boolean;
  signal type_cast_467_inst_req_1 : boolean;
  signal type_cast_467_inst_ack_1 : boolean;
  signal phi_stmt_461_req_1 : boolean;
  signal phi_stmt_461_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "zeropad3D_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  zeropad3D_CP_676_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "zeropad3D_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_CP_676_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= zeropad3D_CP_676_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_CP_676_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  zeropad3D_CP_676: Block -- control-path 
    signal zeropad3D_CP_676_elements: BooleanArray(560 downto 0);
    -- 
  begin -- 
    zeropad3D_CP_676_elements(0) <= zeropad3D_CP_676_start;
    zeropad3D_CP_676_symbol <= zeropad3D_CP_676_elements(553);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	65 
    -- CP-element group 0: 	68 
    -- CP-element group 0: 	29 
    -- CP-element group 0: 	33 
    -- CP-element group 0: 	25 
    -- CP-element group 0: 	39 
    -- CP-element group 0: 	43 
    -- CP-element group 0: 	47 
    -- CP-element group 0: 	51 
    -- CP-element group 0: 	55 
    -- CP-element group 0: 	59 
    -- CP-element group 0: 	62 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	13 
    -- CP-element group 0: 	17 
    -- CP-element group 0: 	21 
    -- CP-element group 0:  members (53) 
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_254_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_224_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_266_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_266_update_start_
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_224_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432__entry__
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_304_update_start_
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_224_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_222/branch_block_stmt_222__entry__
      -- CP-element group 0: 	 branch_block_stmt_222/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_279_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_279_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_241_update_start_
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_241_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_254_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_254_update_start_
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/$entry
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_241_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_266_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_291_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_304_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_304_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_291_update_start_
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_279_update_start_
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_291_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_319_update_start_
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_319_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_319_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_332_update_start_
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_332_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_332_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_344_update_start_
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_344_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_344_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_357_update_start_
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_357_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_357_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_369_update_start_
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_369_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_369_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_382_update_start_
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_382_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_382_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_391_update_start_
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_391_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_391_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_395_update_start_
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_395_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_395_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_399_update_start_
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_399_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_399_Update/cr
      -- 
    cr_833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => type_cast_254_inst_req_1); -- 
    rr_730_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_730_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => RPIPE_zeropad_input_pipe_224_inst_req_0); -- 
    cr_889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => type_cast_279_inst_req_1); -- 
    cr_805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => type_cast_241_inst_req_1); -- 
    cr_861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => type_cast_266_inst_req_1); -- 
    cr_917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => type_cast_291_inst_req_1); -- 
    cr_945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => type_cast_304_inst_req_1); -- 
    cr_987_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_987_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => type_cast_319_inst_req_1); -- 
    cr_1015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => type_cast_332_inst_req_1); -- 
    cr_1043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => type_cast_344_inst_req_1); -- 
    cr_1071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => type_cast_357_inst_req_1); -- 
    cr_1099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => type_cast_369_inst_req_1); -- 
    cr_1127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => type_cast_382_inst_req_1); -- 
    cr_1141_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1141_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => type_cast_391_inst_req_1); -- 
    cr_1155_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1155_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => type_cast_395_inst_req_1); -- 
    cr_1169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => type_cast_399_inst_req_1); -- 
    -- CP-element group 1:  branch  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	499 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	500 
    -- CP-element group 1: 	501 
    -- CP-element group 1:  members (9) 
      -- CP-element group 1: 	 branch_block_stmt_222/if_stmt_1331_eval_test/branch_req
      -- CP-element group 1: 	 branch_block_stmt_222/do_while_stmt_707__exit__
      -- CP-element group 1: 	 branch_block_stmt_222/if_stmt_1331_eval_test/$entry
      -- CP-element group 1: 	 branch_block_stmt_222/if_stmt_1331__entry__
      -- CP-element group 1: 	 branch_block_stmt_222/if_stmt_1331_eval_test/$exit
      -- CP-element group 1: 	 branch_block_stmt_222/if_stmt_1331_dead_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_222/if_stmt_1331_if_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_222/if_stmt_1331_else_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_222/R_ifx_xend304_whilex_xend_taken_1332_place
      -- 
    branch_req_2991_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2991_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(1), ack => if_stmt_1331_branch_req_0); -- 
    zeropad3D_CP_676_elements(1) <= zeropad3D_CP_676_elements(499);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_224_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_224_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_224_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_224_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_224_update_start_
      -- CP-element group 2: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_224_Update/cr
      -- 
    ra_731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_224_inst_ack_0, ack => zeropad3D_CP_676_elements(2)); -- 
    cr_735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(2), ack => RPIPE_zeropad_input_pipe_224_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_224_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_227_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_227_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_227_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_224_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_224_update_completed_
      -- 
    ca_736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_224_inst_ack_1, ack => zeropad3D_CP_676_elements(3)); -- 
    rr_744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(3), ack => RPIPE_zeropad_input_pipe_227_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_227_Update/cr
      -- CP-element group 4: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_227_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_227_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_227_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_227_update_start_
      -- CP-element group 4: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_227_sample_completed_
      -- 
    ra_745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_227_inst_ack_0, ack => zeropad3D_CP_676_elements(4)); -- 
    cr_749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(4), ack => RPIPE_zeropad_input_pipe_227_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_227_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_230_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_227_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_230_Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_230_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_227_update_completed_
      -- 
    ca_750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_227_inst_ack_1, ack => zeropad3D_CP_676_elements(5)); -- 
    rr_758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(5), ack => RPIPE_zeropad_input_pipe_230_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_230_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_230_update_start_
      -- CP-element group 6: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_230_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_230_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_230_Update/cr
      -- CP-element group 6: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_230_Update/$entry
      -- 
    ra_759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_230_inst_ack_0, ack => zeropad3D_CP_676_elements(6)); -- 
    cr_763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(6), ack => RPIPE_zeropad_input_pipe_230_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_233_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_230_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_230_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_230_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_233_Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_233_Sample/$entry
      -- 
    ca_764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_230_inst_ack_1, ack => zeropad3D_CP_676_elements(7)); -- 
    rr_772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(7), ack => RPIPE_zeropad_input_pipe_233_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_233_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_233_update_start_
      -- CP-element group 8: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_233_Update/cr
      -- CP-element group 8: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_233_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_233_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_233_Sample/$exit
      -- 
    ra_773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_233_inst_ack_0, ack => zeropad3D_CP_676_elements(8)); -- 
    cr_777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(8), ack => RPIPE_zeropad_input_pipe_233_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_233_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_233_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_236_Sample/rr
      -- CP-element group 9: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_236_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_233_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_236_sample_start_
      -- 
    ca_778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_233_inst_ack_1, ack => zeropad3D_CP_676_elements(9)); -- 
    rr_786_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_786_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(9), ack => RPIPE_zeropad_input_pipe_236_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_236_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_236_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_236_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_236_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_236_update_start_
      -- CP-element group 10: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_236_sample_completed_
      -- 
    ra_787_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_236_inst_ack_0, ack => zeropad3D_CP_676_elements(10)); -- 
    cr_791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(10), ack => RPIPE_zeropad_input_pipe_236_inst_req_1); -- 
    -- CP-element group 11:  fork  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: 	14 
    -- CP-element group 11:  members (9) 
      -- CP-element group 11: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_236_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_236_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_236_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_241_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_250_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_250_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_241_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_250_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_241_Sample/$entry
      -- 
    ca_792_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_236_inst_ack_1, ack => zeropad3D_CP_676_elements(11)); -- 
    rr_800_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_800_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(11), ack => type_cast_241_inst_req_0); -- 
    rr_814_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_814_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(11), ack => RPIPE_zeropad_input_pipe_250_inst_req_0); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_241_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_241_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_241_Sample/$exit
      -- 
    ra_801_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_241_inst_ack_0, ack => zeropad3D_CP_676_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	0 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	60 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_241_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_241_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_241_Update/$exit
      -- 
    ca_806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_241_inst_ack_1, ack => zeropad3D_CP_676_elements(13)); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	11 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_250_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_250_update_start_
      -- CP-element group 14: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_250_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_250_Update/cr
      -- CP-element group 14: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_250_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_250_Sample/ra
      -- 
    ra_815_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_250_inst_ack_0, ack => zeropad3D_CP_676_elements(14)); -- 
    cr_819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(14), ack => RPIPE_zeropad_input_pipe_250_inst_req_1); -- 
    -- CP-element group 15:  fork  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15: 	18 
    -- CP-element group 15:  members (9) 
      -- CP-element group 15: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_262_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_254_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_254_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_254_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_262_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_250_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_262_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_250_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_250_Update/$exit
      -- 
    ca_820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_250_inst_ack_1, ack => zeropad3D_CP_676_elements(15)); -- 
    rr_828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(15), ack => type_cast_254_inst_req_0); -- 
    rr_842_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_842_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(15), ack => RPIPE_zeropad_input_pipe_262_inst_req_0); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_254_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_254_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_254_sample_completed_
      -- 
    ra_829_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_254_inst_ack_0, ack => zeropad3D_CP_676_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	0 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	60 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_254_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_254_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_254_Update/ca
      -- 
    ca_834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_254_inst_ack_1, ack => zeropad3D_CP_676_elements(17)); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	15 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_262_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_262_Update/cr
      -- CP-element group 18: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_262_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_262_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_262_update_start_
      -- CP-element group 18: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_262_sample_completed_
      -- 
    ra_843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_262_inst_ack_0, ack => zeropad3D_CP_676_elements(18)); -- 
    cr_847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(18), ack => RPIPE_zeropad_input_pipe_262_inst_req_1); -- 
    -- CP-element group 19:  fork  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19: 	22 
    -- CP-element group 19:  members (9) 
      -- CP-element group 19: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_266_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_266_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_266_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_275_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_262_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_262_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_275_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_262_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_275_Sample/$entry
      -- 
    ca_848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_262_inst_ack_1, ack => zeropad3D_CP_676_elements(19)); -- 
    rr_856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(19), ack => type_cast_266_inst_req_0); -- 
    rr_870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(19), ack => RPIPE_zeropad_input_pipe_275_inst_req_0); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_266_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_266_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_266_sample_completed_
      -- 
    ra_857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_266_inst_ack_0, ack => zeropad3D_CP_676_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	0 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	63 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_266_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_266_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_266_Update/ca
      -- 
    ca_862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_266_inst_ack_1, ack => zeropad3D_CP_676_elements(21)); -- 
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	19 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (6) 
      -- CP-element group 22: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_275_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_275_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_275_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_275_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_275_update_start_
      -- CP-element group 22: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_275_Update/cr
      -- 
    ra_871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_275_inst_ack_0, ack => zeropad3D_CP_676_elements(22)); -- 
    cr_875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(22), ack => RPIPE_zeropad_input_pipe_275_inst_req_1); -- 
    -- CP-element group 23:  fork  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: 	26 
    -- CP-element group 23:  members (9) 
      -- CP-element group 23: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_287_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_287_Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_279_Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_279_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_275_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_287_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_275_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_279_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_275_update_completed_
      -- 
    ca_876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_275_inst_ack_1, ack => zeropad3D_CP_676_elements(23)); -- 
    rr_898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(23), ack => RPIPE_zeropad_input_pipe_287_inst_req_0); -- 
    rr_884_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_884_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(23), ack => type_cast_279_inst_req_0); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_279_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_279_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_279_sample_completed_
      -- 
    ra_885_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_279_inst_ack_0, ack => zeropad3D_CP_676_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	0 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	63 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_279_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_279_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_279_Update/ca
      -- 
    ca_890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_279_inst_ack_1, ack => zeropad3D_CP_676_elements(25)); -- 
    -- CP-element group 26:  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	23 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (6) 
      -- CP-element group 26: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_287_update_start_
      -- CP-element group 26: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_287_Update/$entry
      -- CP-element group 26: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_287_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_287_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_287_Update/cr
      -- CP-element group 26: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_287_sample_completed_
      -- 
    ra_899_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_287_inst_ack_0, ack => zeropad3D_CP_676_elements(26)); -- 
    cr_903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(26), ack => RPIPE_zeropad_input_pipe_287_inst_req_1); -- 
    -- CP-element group 27:  fork  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27: 	30 
    -- CP-element group 27:  members (9) 
      -- CP-element group 27: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_291_Sample/rr
      -- CP-element group 27: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_287_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_287_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_287_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_291_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_291_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_300_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_300_Sample/rr
      -- CP-element group 27: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_300_Sample/$entry
      -- 
    ca_904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_287_inst_ack_1, ack => zeropad3D_CP_676_elements(27)); -- 
    rr_912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(27), ack => type_cast_291_inst_req_0); -- 
    rr_926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(27), ack => RPIPE_zeropad_input_pipe_300_inst_req_0); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_291_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_291_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_291_sample_completed_
      -- 
    ra_913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_291_inst_ack_0, ack => zeropad3D_CP_676_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	0 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	66 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_291_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_291_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_291_Update/$exit
      -- 
    ca_918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_291_inst_ack_1, ack => zeropad3D_CP_676_elements(29)); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	27 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_300_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_300_Update/cr
      -- CP-element group 30: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_300_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_300_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_300_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_300_update_start_
      -- 
    ra_927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_300_inst_ack_0, ack => zeropad3D_CP_676_elements(30)); -- 
    cr_931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(30), ack => RPIPE_zeropad_input_pipe_300_inst_req_1); -- 
    -- CP-element group 31:  fork  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31: 	34 
    -- CP-element group 31:  members (9) 
      -- CP-element group 31: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_304_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_304_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_304_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_312_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_312_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_312_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_300_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_300_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_300_update_completed_
      -- 
    ca_932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_300_inst_ack_1, ack => zeropad3D_CP_676_elements(31)); -- 
    rr_940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(31), ack => type_cast_304_inst_req_0); -- 
    rr_954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(31), ack => RPIPE_zeropad_input_pipe_312_inst_req_0); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_304_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_304_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_304_sample_completed_
      -- 
    ra_941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_304_inst_ack_0, ack => zeropad3D_CP_676_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	0 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	66 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_304_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_304_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_304_Update/ca
      -- 
    ca_946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_304_inst_ack_1, ack => zeropad3D_CP_676_elements(33)); -- 
    -- CP-element group 34:  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	31 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (6) 
      -- CP-element group 34: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_312_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_312_update_start_
      -- CP-element group 34: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_312_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_312_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_312_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_312_Sample/ra
      -- 
    ra_955_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_312_inst_ack_0, ack => zeropad3D_CP_676_elements(34)); -- 
    cr_959_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_959_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(34), ack => RPIPE_zeropad_input_pipe_312_inst_req_1); -- 
    -- CP-element group 35:  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (6) 
      -- CP-element group 35: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_312_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_312_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_315_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_315_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_312_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_315_Sample/rr
      -- 
    ca_960_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_312_inst_ack_1, ack => zeropad3D_CP_676_elements(35)); -- 
    rr_968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(35), ack => RPIPE_zeropad_input_pipe_315_inst_req_0); -- 
    -- CP-element group 36:  transition  input  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (6) 
      -- CP-element group 36: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_315_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_315_update_start_
      -- CP-element group 36: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_315_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_315_Sample/ra
      -- CP-element group 36: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_315_Update/$entry
      -- CP-element group 36: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_315_Update/cr
      -- 
    ra_969_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_315_inst_ack_0, ack => zeropad3D_CP_676_elements(36)); -- 
    cr_973_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_973_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(36), ack => RPIPE_zeropad_input_pipe_315_inst_req_1); -- 
    -- CP-element group 37:  fork  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37: 	40 
    -- CP-element group 37:  members (9) 
      -- CP-element group 37: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_315_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_315_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_315_Update/ca
      -- CP-element group 37: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_319_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_319_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_319_Sample/rr
      -- CP-element group 37: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_328_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_328_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_328_Sample/rr
      -- 
    ca_974_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_315_inst_ack_1, ack => zeropad3D_CP_676_elements(37)); -- 
    rr_982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(37), ack => type_cast_319_inst_req_0); -- 
    rr_996_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_996_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(37), ack => RPIPE_zeropad_input_pipe_328_inst_req_0); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_319_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_319_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_319_Sample/ra
      -- 
    ra_983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_319_inst_ack_0, ack => zeropad3D_CP_676_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	0 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	69 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_319_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_319_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_319_Update/ca
      -- 
    ca_988_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_319_inst_ack_1, ack => zeropad3D_CP_676_elements(39)); -- 
    -- CP-element group 40:  transition  input  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	37 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (6) 
      -- CP-element group 40: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_328_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_328_update_start_
      -- CP-element group 40: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_328_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_328_Sample/ra
      -- CP-element group 40: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_328_Update/$entry
      -- CP-element group 40: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_328_Update/cr
      -- 
    ra_997_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_328_inst_ack_0, ack => zeropad3D_CP_676_elements(40)); -- 
    cr_1001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(40), ack => RPIPE_zeropad_input_pipe_328_inst_req_1); -- 
    -- CP-element group 41:  fork  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41: 	44 
    -- CP-element group 41:  members (9) 
      -- CP-element group 41: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_328_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_328_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_328_Update/ca
      -- CP-element group 41: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_332_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_332_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_332_Sample/rr
      -- CP-element group 41: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_340_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_340_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_340_Sample/rr
      -- 
    ca_1002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_328_inst_ack_1, ack => zeropad3D_CP_676_elements(41)); -- 
    rr_1010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(41), ack => type_cast_332_inst_req_0); -- 
    rr_1024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(41), ack => RPIPE_zeropad_input_pipe_340_inst_req_0); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_332_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_332_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_332_Sample/ra
      -- 
    ra_1011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_332_inst_ack_0, ack => zeropad3D_CP_676_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	0 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	69 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_332_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_332_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_332_Update/ca
      -- 
    ca_1016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_332_inst_ack_1, ack => zeropad3D_CP_676_elements(43)); -- 
    -- CP-element group 44:  transition  input  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	41 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (6) 
      -- CP-element group 44: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_340_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_340_update_start_
      -- CP-element group 44: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_340_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_340_Sample/ra
      -- CP-element group 44: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_340_Update/$entry
      -- CP-element group 44: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_340_Update/cr
      -- 
    ra_1025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_340_inst_ack_0, ack => zeropad3D_CP_676_elements(44)); -- 
    cr_1029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(44), ack => RPIPE_zeropad_input_pipe_340_inst_req_1); -- 
    -- CP-element group 45:  fork  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45: 	48 
    -- CP-element group 45:  members (9) 
      -- CP-element group 45: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_340_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_340_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_340_Update/ca
      -- CP-element group 45: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_344_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_344_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_344_Sample/rr
      -- CP-element group 45: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_353_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_353_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_353_Sample/rr
      -- 
    ca_1030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_340_inst_ack_1, ack => zeropad3D_CP_676_elements(45)); -- 
    rr_1038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(45), ack => type_cast_344_inst_req_0); -- 
    rr_1052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(45), ack => RPIPE_zeropad_input_pipe_353_inst_req_0); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_344_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_344_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_344_Sample/ra
      -- 
    ra_1039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_344_inst_ack_0, ack => zeropad3D_CP_676_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	0 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	69 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_344_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_344_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_344_Update/ca
      -- 
    ca_1044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_344_inst_ack_1, ack => zeropad3D_CP_676_elements(47)); -- 
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	45 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (6) 
      -- CP-element group 48: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_353_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_353_update_start_
      -- CP-element group 48: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_353_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_353_Sample/ra
      -- CP-element group 48: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_353_Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_353_Update/cr
      -- 
    ra_1053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_353_inst_ack_0, ack => zeropad3D_CP_676_elements(48)); -- 
    cr_1057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(48), ack => RPIPE_zeropad_input_pipe_353_inst_req_1); -- 
    -- CP-element group 49:  fork  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49: 	52 
    -- CP-element group 49:  members (9) 
      -- CP-element group 49: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_353_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_353_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_353_Update/ca
      -- CP-element group 49: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_357_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_357_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_357_Sample/rr
      -- CP-element group 49: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_365_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_365_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_365_Sample/rr
      -- 
    ca_1058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_353_inst_ack_1, ack => zeropad3D_CP_676_elements(49)); -- 
    rr_1066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(49), ack => type_cast_357_inst_req_0); -- 
    rr_1080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(49), ack => RPIPE_zeropad_input_pipe_365_inst_req_0); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_357_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_357_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_357_Sample/ra
      -- 
    ra_1067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_357_inst_ack_0, ack => zeropad3D_CP_676_elements(50)); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	0 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	69 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_357_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_357_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_357_Update/ca
      -- 
    ca_1072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_357_inst_ack_1, ack => zeropad3D_CP_676_elements(51)); -- 
    -- CP-element group 52:  transition  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	49 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (6) 
      -- CP-element group 52: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_365_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_365_update_start_
      -- CP-element group 52: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_365_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_365_Sample/ra
      -- CP-element group 52: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_365_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_365_Update/cr
      -- 
    ra_1081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_365_inst_ack_0, ack => zeropad3D_CP_676_elements(52)); -- 
    cr_1085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(52), ack => RPIPE_zeropad_input_pipe_365_inst_req_1); -- 
    -- CP-element group 53:  fork  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53: 	56 
    -- CP-element group 53:  members (9) 
      -- CP-element group 53: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_365_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_365_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_365_Update/ca
      -- CP-element group 53: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_369_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_369_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_369_Sample/rr
      -- CP-element group 53: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_378_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_378_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_378_Sample/rr
      -- 
    ca_1086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_365_inst_ack_1, ack => zeropad3D_CP_676_elements(53)); -- 
    rr_1094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(53), ack => type_cast_369_inst_req_0); -- 
    rr_1108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(53), ack => RPIPE_zeropad_input_pipe_378_inst_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_369_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_369_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_369_Sample/ra
      -- 
    ra_1095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_369_inst_ack_0, ack => zeropad3D_CP_676_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	0 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	69 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_369_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_369_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_369_Update/ca
      -- 
    ca_1100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_369_inst_ack_1, ack => zeropad3D_CP_676_elements(55)); -- 
    -- CP-element group 56:  transition  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	53 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (6) 
      -- CP-element group 56: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_378_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_378_update_start_
      -- CP-element group 56: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_378_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_378_Sample/ra
      -- CP-element group 56: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_378_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_378_Update/cr
      -- 
    ra_1109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_378_inst_ack_0, ack => zeropad3D_CP_676_elements(56)); -- 
    cr_1113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(56), ack => RPIPE_zeropad_input_pipe_378_inst_req_1); -- 
    -- CP-element group 57:  transition  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (6) 
      -- CP-element group 57: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_378_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_378_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/RPIPE_zeropad_input_pipe_378_Update/ca
      -- CP-element group 57: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_382_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_382_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_382_Sample/rr
      -- 
    ca_1114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_378_inst_ack_1, ack => zeropad3D_CP_676_elements(57)); -- 
    rr_1122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(57), ack => type_cast_382_inst_req_0); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_382_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_382_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_382_Sample/ra
      -- 
    ra_1123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_382_inst_ack_0, ack => zeropad3D_CP_676_elements(58)); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	0 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	69 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_382_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_382_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_382_Update/ca
      -- 
    ca_1128_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_382_inst_ack_1, ack => zeropad3D_CP_676_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	13 
    -- CP-element group 60: 	17 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_391_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_391_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_391_Sample/rr
      -- 
    rr_1136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(60), ack => type_cast_391_inst_req_0); -- 
    zeropad3D_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(13) & zeropad3D_CP_676_elements(17);
      gj_zeropad3D_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_391_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_391_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_391_Sample/ra
      -- 
    ra_1137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_391_inst_ack_0, ack => zeropad3D_CP_676_elements(61)); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	0 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	69 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_391_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_391_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_391_Update/ca
      -- 
    ca_1142_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_391_inst_ack_1, ack => zeropad3D_CP_676_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	25 
    -- CP-element group 63: 	21 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_395_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_395_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_395_Sample/rr
      -- 
    rr_1150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(63), ack => type_cast_395_inst_req_0); -- 
    zeropad3D_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(25) & zeropad3D_CP_676_elements(21);
      gj_zeropad3D_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_395_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_395_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_395_Sample/ra
      -- 
    ra_1151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_395_inst_ack_0, ack => zeropad3D_CP_676_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	0 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	69 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_395_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_395_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_395_Update/ca
      -- 
    ca_1156_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_395_inst_ack_1, ack => zeropad3D_CP_676_elements(65)); -- 
    -- CP-element group 66:  join  transition  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	29 
    -- CP-element group 66: 	33 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_399_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_399_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_399_Sample/rr
      -- 
    rr_1164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(66), ack => type_cast_399_inst_req_0); -- 
    zeropad3D_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(29) & zeropad3D_CP_676_elements(33);
      gj_zeropad3D_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_399_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_399_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_399_Sample/ra
      -- 
    ra_1165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_399_inst_ack_0, ack => zeropad3D_CP_676_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	0 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_399_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_399_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/type_cast_399_Update/ca
      -- 
    ca_1170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_399_inst_ack_1, ack => zeropad3D_CP_676_elements(68)); -- 
    -- CP-element group 69:  branch  join  transition  place  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	65 
    -- CP-element group 69: 	68 
    -- CP-element group 69: 	39 
    -- CP-element group 69: 	43 
    -- CP-element group 69: 	47 
    -- CP-element group 69: 	51 
    -- CP-element group 69: 	55 
    -- CP-element group 69: 	59 
    -- CP-element group 69: 	62 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (10) 
      -- CP-element group 69: 	 branch_block_stmt_222/if_stmt_433__entry__
      -- CP-element group 69: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432__exit__
      -- CP-element group 69: 	 branch_block_stmt_222/assign_stmt_225_to_assign_stmt_432/$exit
      -- CP-element group 69: 	 branch_block_stmt_222/if_stmt_433_dead_link/$entry
      -- CP-element group 69: 	 branch_block_stmt_222/if_stmt_433_eval_test/$entry
      -- CP-element group 69: 	 branch_block_stmt_222/if_stmt_433_eval_test/$exit
      -- CP-element group 69: 	 branch_block_stmt_222/if_stmt_433_eval_test/branch_req
      -- CP-element group 69: 	 branch_block_stmt_222/R_cmp390_434_place
      -- CP-element group 69: 	 branch_block_stmt_222/if_stmt_433_if_link/$entry
      -- CP-element group 69: 	 branch_block_stmt_222/if_stmt_433_else_link/$entry
      -- 
    branch_req_1178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(69), ack => if_stmt_433_branch_req_0); -- 
    zeropad3D_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(65) & zeropad3D_CP_676_elements(68) & zeropad3D_CP_676_elements(39) & zeropad3D_CP_676_elements(43) & zeropad3D_CP_676_elements(47) & zeropad3D_CP_676_elements(51) & zeropad3D_CP_676_elements(55) & zeropad3D_CP_676_elements(59) & zeropad3D_CP_676_elements(62);
      gj_zeropad3D_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  merge  transition  place  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	554 
    -- CP-element group 70:  members (18) 
      -- CP-element group 70: 	 branch_block_stmt_222/assign_stmt_445_to_assign_stmt_458__entry__
      -- CP-element group 70: 	 branch_block_stmt_222/merge_stmt_439__exit__
      -- CP-element group 70: 	 branch_block_stmt_222/bbx_xnph_forx_xbody
      -- CP-element group 70: 	 branch_block_stmt_222/assign_stmt_445_to_assign_stmt_458__exit__
      -- CP-element group 70: 	 branch_block_stmt_222/if_stmt_433_if_link/$exit
      -- CP-element group 70: 	 branch_block_stmt_222/if_stmt_433_if_link/if_choice_transition
      -- CP-element group 70: 	 branch_block_stmt_222/entry_bbx_xnph
      -- CP-element group 70: 	 branch_block_stmt_222/assign_stmt_445_to_assign_stmt_458/$entry
      -- CP-element group 70: 	 branch_block_stmt_222/assign_stmt_445_to_assign_stmt_458/$exit
      -- CP-element group 70: 	 branch_block_stmt_222/entry_bbx_xnph_PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_222/entry_bbx_xnph_PhiReq/$exit
      -- CP-element group 70: 	 branch_block_stmt_222/merge_stmt_439_PhiReqMerge
      -- CP-element group 70: 	 branch_block_stmt_222/merge_stmt_439_PhiAck/$entry
      -- CP-element group 70: 	 branch_block_stmt_222/merge_stmt_439_PhiAck/$exit
      -- CP-element group 70: 	 branch_block_stmt_222/merge_stmt_439_PhiAck/dummy
      -- CP-element group 70: 	 branch_block_stmt_222/bbx_xnph_forx_xbody_PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_222/bbx_xnph_forx_xbody_PhiReq/phi_stmt_461/$entry
      -- CP-element group 70: 	 branch_block_stmt_222/bbx_xnph_forx_xbody_PhiReq/phi_stmt_461/phi_stmt_461_sources/$entry
      -- 
    if_choice_transition_1183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_433_branch_ack_1, ack => zeropad3D_CP_676_elements(70)); -- 
    -- CP-element group 71:  transition  place  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	560 
    -- CP-element group 71:  members (5) 
      -- CP-element group 71: 	 branch_block_stmt_222/if_stmt_433_else_link/$exit
      -- CP-element group 71: 	 branch_block_stmt_222/if_stmt_433_else_link/else_choice_transition
      -- CP-element group 71: 	 branch_block_stmt_222/entry_forx_xend
      -- CP-element group 71: 	 branch_block_stmt_222/entry_forx_xend_PhiReq/$entry
      -- CP-element group 71: 	 branch_block_stmt_222/entry_forx_xend_PhiReq/$exit
      -- 
    else_choice_transition_1187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_433_branch_ack_0, ack => zeropad3D_CP_676_elements(71)); -- 
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	559 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	111 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/array_obj_ref_473_final_index_sum_regn_sample_complete
      -- CP-element group 72: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/array_obj_ref_473_final_index_sum_regn_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/array_obj_ref_473_final_index_sum_regn_Sample/ack
      -- 
    ack_1221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_473_index_offset_ack_0, ack => zeropad3D_CP_676_elements(72)); -- 
    -- CP-element group 73:  transition  input  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	559 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (11) 
      -- CP-element group 73: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/addr_of_474_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/array_obj_ref_473_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/array_obj_ref_473_offset_calculated
      -- CP-element group 73: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/array_obj_ref_473_final_index_sum_regn_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/array_obj_ref_473_final_index_sum_regn_Update/ack
      -- CP-element group 73: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/array_obj_ref_473_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/array_obj_ref_473_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/array_obj_ref_473_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/array_obj_ref_473_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/addr_of_474_request/$entry
      -- CP-element group 73: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/addr_of_474_request/req
      -- 
    ack_1226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_473_index_offset_ack_1, ack => zeropad3D_CP_676_elements(73)); -- 
    req_1235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(73), ack => addr_of_474_final_reg_req_0); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/addr_of_474_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/addr_of_474_request/$exit
      -- CP-element group 74: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/addr_of_474_request/ack
      -- 
    ack_1236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_474_final_reg_ack_0, ack => zeropad3D_CP_676_elements(74)); -- 
    -- CP-element group 75:  fork  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	559 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	108 
    -- CP-element group 75:  members (19) 
      -- CP-element group 75: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/ptr_deref_610_word_addrgen/root_register_ack
      -- CP-element group 75: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/ptr_deref_610_base_plus_offset/$exit
      -- CP-element group 75: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/ptr_deref_610_word_addrgen/root_register_req
      -- CP-element group 75: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/ptr_deref_610_base_plus_offset/sum_rename_ack
      -- CP-element group 75: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/ptr_deref_610_word_addrgen/$entry
      -- CP-element group 75: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/ptr_deref_610_word_addrgen/$exit
      -- CP-element group 75: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/ptr_deref_610_base_plus_offset/sum_rename_req
      -- CP-element group 75: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/ptr_deref_610_base_plus_offset/$entry
      -- CP-element group 75: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/ptr_deref_610_base_addr_resize/base_resize_ack
      -- CP-element group 75: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/addr_of_474_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/ptr_deref_610_base_addr_resize/base_resize_req
      -- CP-element group 75: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/ptr_deref_610_base_addr_resize/$exit
      -- CP-element group 75: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/addr_of_474_complete/$exit
      -- CP-element group 75: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/addr_of_474_complete/ack
      -- CP-element group 75: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/ptr_deref_610_base_address_calculated
      -- CP-element group 75: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/ptr_deref_610_word_address_calculated
      -- CP-element group 75: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/ptr_deref_610_root_address_calculated
      -- CP-element group 75: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/ptr_deref_610_base_address_resized
      -- CP-element group 75: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/ptr_deref_610_base_addr_resize/$entry
      -- 
    ack_1241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_474_final_reg_ack_1, ack => zeropad3D_CP_676_elements(75)); -- 
    -- CP-element group 76:  transition  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	559 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (6) 
      -- CP-element group 76: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_477_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_477_update_start_
      -- CP-element group 76: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_477_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_477_Sample/ra
      -- CP-element group 76: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_477_Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_477_Update/cr
      -- 
    ra_1250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_477_inst_ack_0, ack => zeropad3D_CP_676_elements(76)); -- 
    cr_1254_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1254_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(76), ack => RPIPE_zeropad_input_pipe_477_inst_req_1); -- 
    -- CP-element group 77:  fork  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	80 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (9) 
      -- CP-element group 77: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_477_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_477_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_477_Update/ca
      -- CP-element group 77: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_481_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_481_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_481_Sample/rr
      -- CP-element group 77: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_490_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_490_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_490_Sample/rr
      -- 
    ca_1255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_477_inst_ack_1, ack => zeropad3D_CP_676_elements(77)); -- 
    rr_1277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(77), ack => RPIPE_zeropad_input_pipe_490_inst_req_0); -- 
    rr_1263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(77), ack => type_cast_481_inst_req_0); -- 
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_481_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_481_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_481_Sample/ra
      -- 
    ra_1264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_481_inst_ack_0, ack => zeropad3D_CP_676_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	559 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	108 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_481_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_481_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_481_Update/ca
      -- 
    ca_1269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_481_inst_ack_1, ack => zeropad3D_CP_676_elements(79)); -- 
    -- CP-element group 80:  transition  input  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	77 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (6) 
      -- CP-element group 80: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_490_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_490_update_start_
      -- CP-element group 80: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_490_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_490_Sample/ra
      -- CP-element group 80: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_490_Update/$entry
      -- CP-element group 80: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_490_Update/cr
      -- 
    ra_1278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_490_inst_ack_0, ack => zeropad3D_CP_676_elements(80)); -- 
    cr_1282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(80), ack => RPIPE_zeropad_input_pipe_490_inst_req_1); -- 
    -- CP-element group 81:  fork  transition  input  output  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	84 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (9) 
      -- CP-element group 81: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_490_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_490_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_490_Update/ca
      -- CP-element group 81: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_494_sample_start_
      -- CP-element group 81: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_494_Sample/$entry
      -- CP-element group 81: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_494_Sample/rr
      -- CP-element group 81: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_508_sample_start_
      -- CP-element group 81: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_508_Sample/$entry
      -- CP-element group 81: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_508_Sample/rr
      -- 
    ca_1283_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_490_inst_ack_1, ack => zeropad3D_CP_676_elements(81)); -- 
    rr_1291_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1291_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(81), ack => type_cast_494_inst_req_0); -- 
    rr_1305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(81), ack => RPIPE_zeropad_input_pipe_508_inst_req_0); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_494_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_494_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_494_Sample/ra
      -- 
    ra_1292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_494_inst_ack_0, ack => zeropad3D_CP_676_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	559 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	108 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_494_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_494_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_494_Update/ca
      -- 
    ca_1297_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_494_inst_ack_1, ack => zeropad3D_CP_676_elements(83)); -- 
    -- CP-element group 84:  transition  input  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	81 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (6) 
      -- CP-element group 84: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_508_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_508_update_start_
      -- CP-element group 84: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_508_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_508_Sample/ra
      -- CP-element group 84: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_508_Update/$entry
      -- CP-element group 84: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_508_Update/cr
      -- 
    ra_1306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_508_inst_ack_0, ack => zeropad3D_CP_676_elements(84)); -- 
    cr_1310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(84), ack => RPIPE_zeropad_input_pipe_508_inst_req_1); -- 
    -- CP-element group 85:  fork  transition  input  output  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	88 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (9) 
      -- CP-element group 85: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_508_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_508_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_508_Update/ca
      -- CP-element group 85: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_512_sample_start_
      -- CP-element group 85: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_512_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_512_Sample/rr
      -- CP-element group 85: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_526_sample_start_
      -- CP-element group 85: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_526_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_526_Sample/rr
      -- 
    ca_1311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_508_inst_ack_1, ack => zeropad3D_CP_676_elements(85)); -- 
    rr_1333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(85), ack => RPIPE_zeropad_input_pipe_526_inst_req_0); -- 
    rr_1319_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1319_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(85), ack => type_cast_512_inst_req_0); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_512_sample_completed_
      -- CP-element group 86: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_512_Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_512_Sample/ra
      -- 
    ra_1320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_512_inst_ack_0, ack => zeropad3D_CP_676_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	559 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	108 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_512_update_completed_
      -- CP-element group 87: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_512_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_512_Update/ca
      -- 
    ca_1325_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_512_inst_ack_1, ack => zeropad3D_CP_676_elements(87)); -- 
    -- CP-element group 88:  transition  input  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	85 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (6) 
      -- CP-element group 88: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_526_sample_completed_
      -- CP-element group 88: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_526_update_start_
      -- CP-element group 88: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_526_Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_526_Sample/ra
      -- CP-element group 88: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_526_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_526_Update/cr
      -- 
    ra_1334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_526_inst_ack_0, ack => zeropad3D_CP_676_elements(88)); -- 
    cr_1338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(88), ack => RPIPE_zeropad_input_pipe_526_inst_req_1); -- 
    -- CP-element group 89:  fork  transition  input  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89: 	92 
    -- CP-element group 89:  members (9) 
      -- CP-element group 89: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_526_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_526_Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_526_Update/ca
      -- CP-element group 89: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_530_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_530_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_530_Sample/rr
      -- CP-element group 89: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_544_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_544_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_544_Sample/rr
      -- 
    ca_1339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_526_inst_ack_1, ack => zeropad3D_CP_676_elements(89)); -- 
    rr_1347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(89), ack => type_cast_530_inst_req_0); -- 
    rr_1361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(89), ack => RPIPE_zeropad_input_pipe_544_inst_req_0); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_530_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_530_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_530_Sample/ra
      -- 
    ra_1348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_530_inst_ack_0, ack => zeropad3D_CP_676_elements(90)); -- 
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	559 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	108 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_530_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_530_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_530_Update/ca
      -- 
    ca_1353_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_530_inst_ack_1, ack => zeropad3D_CP_676_elements(91)); -- 
    -- CP-element group 92:  transition  input  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	89 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92:  members (6) 
      -- CP-element group 92: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_544_sample_completed_
      -- CP-element group 92: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_544_update_start_
      -- CP-element group 92: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_544_Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_544_Sample/ra
      -- CP-element group 92: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_544_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_544_Update/cr
      -- 
    ra_1362_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_544_inst_ack_0, ack => zeropad3D_CP_676_elements(92)); -- 
    cr_1366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(92), ack => RPIPE_zeropad_input_pipe_544_inst_req_1); -- 
    -- CP-element group 93:  fork  transition  input  output  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93: 	96 
    -- CP-element group 93:  members (9) 
      -- CP-element group 93: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_544_update_completed_
      -- CP-element group 93: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_544_Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_544_Update/ca
      -- CP-element group 93: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_548_sample_start_
      -- CP-element group 93: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_548_Sample/$entry
      -- CP-element group 93: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_548_Sample/rr
      -- CP-element group 93: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_562_sample_start_
      -- CP-element group 93: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_562_Sample/$entry
      -- CP-element group 93: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_562_Sample/rr
      -- 
    ca_1367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_544_inst_ack_1, ack => zeropad3D_CP_676_elements(93)); -- 
    rr_1375_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1375_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(93), ack => type_cast_548_inst_req_0); -- 
    rr_1389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(93), ack => RPIPE_zeropad_input_pipe_562_inst_req_0); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_548_sample_completed_
      -- CP-element group 94: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_548_Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_548_Sample/ra
      -- 
    ra_1376_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_548_inst_ack_0, ack => zeropad3D_CP_676_elements(94)); -- 
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	559 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	108 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_548_update_completed_
      -- CP-element group 95: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_548_Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_548_Update/ca
      -- 
    ca_1381_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_548_inst_ack_1, ack => zeropad3D_CP_676_elements(95)); -- 
    -- CP-element group 96:  transition  input  output  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	93 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (6) 
      -- CP-element group 96: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_562_sample_completed_
      -- CP-element group 96: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_562_update_start_
      -- CP-element group 96: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_562_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_562_Sample/ra
      -- CP-element group 96: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_562_Update/$entry
      -- CP-element group 96: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_562_Update/cr
      -- 
    ra_1390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_562_inst_ack_0, ack => zeropad3D_CP_676_elements(96)); -- 
    cr_1394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(96), ack => RPIPE_zeropad_input_pipe_562_inst_req_1); -- 
    -- CP-element group 97:  fork  transition  input  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97: 	100 
    -- CP-element group 97:  members (9) 
      -- CP-element group 97: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_562_update_completed_
      -- CP-element group 97: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_562_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_562_Update/ca
      -- CP-element group 97: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_566_sample_start_
      -- CP-element group 97: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_566_Sample/$entry
      -- CP-element group 97: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_566_Sample/rr
      -- CP-element group 97: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_580_sample_start_
      -- CP-element group 97: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_580_Sample/$entry
      -- CP-element group 97: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_580_Sample/rr
      -- 
    ca_1395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_562_inst_ack_1, ack => zeropad3D_CP_676_elements(97)); -- 
    rr_1403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(97), ack => type_cast_566_inst_req_0); -- 
    rr_1417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(97), ack => RPIPE_zeropad_input_pipe_580_inst_req_0); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_566_sample_completed_
      -- CP-element group 98: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_566_Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_566_Sample/ra
      -- 
    ra_1404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_566_inst_ack_0, ack => zeropad3D_CP_676_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	559 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	108 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_566_update_completed_
      -- CP-element group 99: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_566_Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_566_Update/ca
      -- 
    ca_1409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_566_inst_ack_1, ack => zeropad3D_CP_676_elements(99)); -- 
    -- CP-element group 100:  transition  input  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	97 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100:  members (6) 
      -- CP-element group 100: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_580_sample_completed_
      -- CP-element group 100: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_580_update_start_
      -- CP-element group 100: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_580_Sample/$exit
      -- CP-element group 100: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_580_Sample/ra
      -- CP-element group 100: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_580_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_580_Update/cr
      -- 
    ra_1418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_580_inst_ack_0, ack => zeropad3D_CP_676_elements(100)); -- 
    cr_1422_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1422_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(100), ack => RPIPE_zeropad_input_pipe_580_inst_req_1); -- 
    -- CP-element group 101:  fork  transition  input  output  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	102 
    -- CP-element group 101: 	104 
    -- CP-element group 101:  members (9) 
      -- CP-element group 101: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_580_update_completed_
      -- CP-element group 101: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_580_Update/$exit
      -- CP-element group 101: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_580_Update/ca
      -- CP-element group 101: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_584_sample_start_
      -- CP-element group 101: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_584_Sample/$entry
      -- CP-element group 101: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_584_Sample/rr
      -- CP-element group 101: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_598_sample_start_
      -- CP-element group 101: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_598_Sample/$entry
      -- CP-element group 101: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_598_Sample/rr
      -- 
    ca_1423_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_580_inst_ack_1, ack => zeropad3D_CP_676_elements(101)); -- 
    rr_1431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(101), ack => type_cast_584_inst_req_0); -- 
    rr_1445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(101), ack => RPIPE_zeropad_input_pipe_598_inst_req_0); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	101 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_584_sample_completed_
      -- CP-element group 102: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_584_Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_584_Sample/ra
      -- 
    ra_1432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_584_inst_ack_0, ack => zeropad3D_CP_676_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	559 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	108 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_584_update_completed_
      -- CP-element group 103: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_584_Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_584_Update/ca
      -- 
    ca_1437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_584_inst_ack_1, ack => zeropad3D_CP_676_elements(103)); -- 
    -- CP-element group 104:  transition  input  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	101 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (6) 
      -- CP-element group 104: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_598_sample_completed_
      -- CP-element group 104: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_598_update_start_
      -- CP-element group 104: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_598_Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_598_Sample/ra
      -- CP-element group 104: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_598_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_598_Update/cr
      -- 
    ra_1446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_598_inst_ack_0, ack => zeropad3D_CP_676_elements(104)); -- 
    cr_1450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(104), ack => RPIPE_zeropad_input_pipe_598_inst_req_1); -- 
    -- CP-element group 105:  transition  input  output  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	106 
    -- CP-element group 105:  members (6) 
      -- CP-element group 105: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_598_update_completed_
      -- CP-element group 105: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_598_Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_598_Update/ca
      -- CP-element group 105: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_602_sample_start_
      -- CP-element group 105: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_602_Sample/$entry
      -- CP-element group 105: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_602_Sample/rr
      -- 
    ca_1451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_598_inst_ack_1, ack => zeropad3D_CP_676_elements(105)); -- 
    rr_1459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(105), ack => type_cast_602_inst_req_0); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	105 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_602_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_602_Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_602_Sample/ra
      -- 
    ra_1460_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_602_inst_ack_0, ack => zeropad3D_CP_676_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	559 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_602_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_602_Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_602_Update/ca
      -- 
    ca_1465_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_602_inst_ack_1, ack => zeropad3D_CP_676_elements(107)); -- 
    -- CP-element group 108:  join  transition  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	79 
    -- CP-element group 108: 	91 
    -- CP-element group 108: 	95 
    -- CP-element group 108: 	87 
    -- CP-element group 108: 	83 
    -- CP-element group 108: 	75 
    -- CP-element group 108: 	99 
    -- CP-element group 108: 	103 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (9) 
      -- CP-element group 108: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/ptr_deref_610_Sample/ptr_deref_610_Split/$exit
      -- CP-element group 108: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/ptr_deref_610_Sample/ptr_deref_610_Split/split_req
      -- CP-element group 108: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/ptr_deref_610_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/ptr_deref_610_Sample/ptr_deref_610_Split/$entry
      -- CP-element group 108: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/ptr_deref_610_Sample/ptr_deref_610_Split/split_ack
      -- CP-element group 108: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/ptr_deref_610_Sample/word_access_start/word_0/rr
      -- CP-element group 108: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/ptr_deref_610_Sample/word_access_start/word_0/$entry
      -- CP-element group 108: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/ptr_deref_610_Sample/word_access_start/$entry
      -- CP-element group 108: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/ptr_deref_610_sample_start_
      -- 
    rr_1503_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1503_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(108), ack => ptr_deref_610_store_0_req_0); -- 
    zeropad3D_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(79) & zeropad3D_CP_676_elements(91) & zeropad3D_CP_676_elements(95) & zeropad3D_CP_676_elements(87) & zeropad3D_CP_676_elements(83) & zeropad3D_CP_676_elements(75) & zeropad3D_CP_676_elements(99) & zeropad3D_CP_676_elements(103) & zeropad3D_CP_676_elements(107);
      gj_zeropad3D_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (5) 
      -- CP-element group 109: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/ptr_deref_610_Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/ptr_deref_610_Sample/word_access_start/word_0/ra
      -- CP-element group 109: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/ptr_deref_610_Sample/word_access_start/word_0/$exit
      -- CP-element group 109: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/ptr_deref_610_Sample/word_access_start/$exit
      -- CP-element group 109: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/ptr_deref_610_sample_completed_
      -- 
    ra_1504_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_610_store_0_ack_0, ack => zeropad3D_CP_676_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	559 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (5) 
      -- CP-element group 110: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/ptr_deref_610_Update/word_access_complete/word_0/ca
      -- CP-element group 110: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/ptr_deref_610_Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/ptr_deref_610_Update/word_access_complete/$exit
      -- CP-element group 110: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/ptr_deref_610_Update/word_access_complete/word_0/$exit
      -- CP-element group 110: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/ptr_deref_610_update_completed_
      -- 
    ca_1515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_610_store_0_ack_1, ack => zeropad3D_CP_676_elements(110)); -- 
    -- CP-element group 111:  branch  join  transition  place  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	72 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111: 	113 
    -- CP-element group 111:  members (10) 
      -- CP-element group 111: 	 branch_block_stmt_222/if_stmt_624_dead_link/$entry
      -- CP-element group 111: 	 branch_block_stmt_222/if_stmt_624_eval_test/$entry
      -- CP-element group 111: 	 branch_block_stmt_222/if_stmt_624__entry__
      -- CP-element group 111: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623__exit__
      -- CP-element group 111: 	 branch_block_stmt_222/R_exitcond3_625_place
      -- CP-element group 111: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/$exit
      -- CP-element group 111: 	 branch_block_stmt_222/if_stmt_624_else_link/$entry
      -- CP-element group 111: 	 branch_block_stmt_222/if_stmt_624_if_link/$entry
      -- CP-element group 111: 	 branch_block_stmt_222/if_stmt_624_eval_test/branch_req
      -- CP-element group 111: 	 branch_block_stmt_222/if_stmt_624_eval_test/$exit
      -- 
    branch_req_1523_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1523_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(111), ack => if_stmt_624_branch_req_0); -- 
    zeropad3D_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(72) & zeropad3D_CP_676_elements(110);
      gj_zeropad3D_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  merge  transition  place  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	560 
    -- CP-element group 112:  members (13) 
      -- CP-element group 112: 	 branch_block_stmt_222/forx_xendx_xloopexit_forx_xend
      -- CP-element group 112: 	 branch_block_stmt_222/merge_stmt_630__exit__
      -- CP-element group 112: 	 branch_block_stmt_222/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 112: 	 branch_block_stmt_222/if_stmt_624_if_link/if_choice_transition
      -- CP-element group 112: 	 branch_block_stmt_222/if_stmt_624_if_link/$exit
      -- CP-element group 112: 	 branch_block_stmt_222/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 112: 	 branch_block_stmt_222/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 112: 	 branch_block_stmt_222/merge_stmt_630_PhiReqMerge
      -- CP-element group 112: 	 branch_block_stmt_222/merge_stmt_630_PhiAck/$entry
      -- CP-element group 112: 	 branch_block_stmt_222/merge_stmt_630_PhiAck/$exit
      -- CP-element group 112: 	 branch_block_stmt_222/merge_stmt_630_PhiAck/dummy
      -- CP-element group 112: 	 branch_block_stmt_222/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 112: 	 branch_block_stmt_222/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_1528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_624_branch_ack_1, ack => zeropad3D_CP_676_elements(112)); -- 
    -- CP-element group 113:  fork  transition  place  input  output  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	111 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	555 
    -- CP-element group 113: 	556 
    -- CP-element group 113:  members (12) 
      -- CP-element group 113: 	 branch_block_stmt_222/forx_xbody_forx_xbody
      -- CP-element group 113: 	 branch_block_stmt_222/if_stmt_624_else_link/else_choice_transition
      -- CP-element group 113: 	 branch_block_stmt_222/if_stmt_624_else_link/$exit
      -- CP-element group 113: 	 branch_block_stmt_222/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 113: 	 branch_block_stmt_222/forx_xbody_forx_xbody_PhiReq/phi_stmt_461/$entry
      -- CP-element group 113: 	 branch_block_stmt_222/forx_xbody_forx_xbody_PhiReq/phi_stmt_461/phi_stmt_461_sources/$entry
      -- CP-element group 113: 	 branch_block_stmt_222/forx_xbody_forx_xbody_PhiReq/phi_stmt_461/phi_stmt_461_sources/type_cast_467/$entry
      -- CP-element group 113: 	 branch_block_stmt_222/forx_xbody_forx_xbody_PhiReq/phi_stmt_461/phi_stmt_461_sources/type_cast_467/SplitProtocol/$entry
      -- CP-element group 113: 	 branch_block_stmt_222/forx_xbody_forx_xbody_PhiReq/phi_stmt_461/phi_stmt_461_sources/type_cast_467/SplitProtocol/Sample/$entry
      -- CP-element group 113: 	 branch_block_stmt_222/forx_xbody_forx_xbody_PhiReq/phi_stmt_461/phi_stmt_461_sources/type_cast_467/SplitProtocol/Sample/rr
      -- CP-element group 113: 	 branch_block_stmt_222/forx_xbody_forx_xbody_PhiReq/phi_stmt_461/phi_stmt_461_sources/type_cast_467/SplitProtocol/Update/$entry
      -- CP-element group 113: 	 branch_block_stmt_222/forx_xbody_forx_xbody_PhiReq/phi_stmt_461/phi_stmt_461_sources/type_cast_467/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_624_branch_ack_0, ack => zeropad3D_CP_676_elements(113)); -- 
    rr_3360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(113), ack => type_cast_467_inst_req_0); -- 
    cr_3365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(113), ack => type_cast_467_inst_req_1); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	560 
    -- CP-element group 114: successors 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/call_stmt_635_Sample/cra
      -- CP-element group 114: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/call_stmt_635_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/call_stmt_635_sample_completed_
      -- 
    cra_1546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_635_call_ack_0, ack => zeropad3D_CP_676_elements(114)); -- 
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	560 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	126 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/call_stmt_635_Update/cca
      -- CP-element group 115: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/call_stmt_635_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/call_stmt_635_update_completed_
      -- 
    cca_1551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_635_call_ack_1, ack => zeropad3D_CP_676_elements(115)); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	560 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_645_sample_completed_
      -- CP-element group 116: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_645_Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_645_Sample/ra
      -- 
    ra_1560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_645_inst_ack_0, ack => zeropad3D_CP_676_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	560 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	126 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_645_Update/ca
      -- CP-element group 117: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_645_Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_645_update_completed_
      -- 
    ca_1565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_645_inst_ack_1, ack => zeropad3D_CP_676_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	560 
    -- CP-element group 118: successors 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_649_Sample/$exit
      -- CP-element group 118: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_649_Sample/ra
      -- CP-element group 118: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_649_sample_completed_
      -- 
    ra_1574_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_649_inst_ack_0, ack => zeropad3D_CP_676_elements(118)); -- 
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	560 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	126 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_649_update_completed_
      -- CP-element group 119: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_649_Update/$exit
      -- CP-element group 119: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_649_Update/ca
      -- 
    ca_1579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_649_inst_ack_1, ack => zeropad3D_CP_676_elements(119)); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	560 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_653_Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_653_sample_completed_
      -- CP-element group 120: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_653_Sample/ra
      -- 
    ra_1588_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_653_inst_ack_0, ack => zeropad3D_CP_676_elements(120)); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	560 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	126 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_653_update_completed_
      -- CP-element group 121: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_653_Update/$exit
      -- CP-element group 121: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_653_Update/ca
      -- 
    ca_1593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_653_inst_ack_1, ack => zeropad3D_CP_676_elements(121)); -- 
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	560 
    -- CP-element group 122: successors 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_668_sample_completed_
      -- CP-element group 122: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_668_Sample/ra
      -- CP-element group 122: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_668_Sample/$exit
      -- 
    ra_1602_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_668_inst_ack_0, ack => zeropad3D_CP_676_elements(122)); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	560 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	126 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_668_Update/ca
      -- CP-element group 123: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_668_Update/$exit
      -- CP-element group 123: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_668_update_completed_
      -- 
    ca_1607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_668_inst_ack_1, ack => zeropad3D_CP_676_elements(123)); -- 
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	560 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_677_Sample/ra
      -- CP-element group 124: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_677_Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_677_sample_completed_
      -- 
    ra_1616_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_677_inst_ack_0, ack => zeropad3D_CP_676_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	560 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	126 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_677_Update/ca
      -- CP-element group 125: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_677_Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_677_update_completed_
      -- 
    ca_1621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_677_inst_ack_1, ack => zeropad3D_CP_676_elements(125)); -- 
    -- CP-element group 126:  join  transition  place  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	115 
    -- CP-element group 126: 	117 
    -- CP-element group 126: 	119 
    -- CP-element group 126: 	121 
    -- CP-element group 126: 	123 
    -- CP-element group 126: 	125 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (10) 
      -- CP-element group 126: 	 branch_block_stmt_222/do_while_stmt_707__entry__
      -- CP-element group 126: 	 branch_block_stmt_222/merge_stmt_690__exit__
      -- CP-element group 126: 	 branch_block_stmt_222/forx_xend_whilex_xbody
      -- CP-element group 126: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688__exit__
      -- CP-element group 126: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/$exit
      -- CP-element group 126: 	 branch_block_stmt_222/forx_xend_whilex_xbody_PhiReq/$entry
      -- CP-element group 126: 	 branch_block_stmt_222/forx_xend_whilex_xbody_PhiReq/$exit
      -- CP-element group 126: 	 branch_block_stmt_222/merge_stmt_690_PhiReqMerge
      -- CP-element group 126: 	 branch_block_stmt_222/merge_stmt_690_PhiAck/$entry
      -- CP-element group 126: 	 branch_block_stmt_222/merge_stmt_690_PhiAck/$exit
      -- 
    zeropad3D_cp_element_group_126: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_126"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(115) & zeropad3D_CP_676_elements(117) & zeropad3D_CP_676_elements(119) & zeropad3D_CP_676_elements(121) & zeropad3D_CP_676_elements(123) & zeropad3D_CP_676_elements(125);
      gj_zeropad3D_cp_element_group_126 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(126), clk => clk, reset => reset); --
    end block;
    -- CP-element group 127:  transition  place  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	133 
    -- CP-element group 127:  members (2) 
      -- CP-element group 127: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707__entry__
      -- CP-element group 127: 	 branch_block_stmt_222/do_while_stmt_707/$entry
      -- 
    zeropad3D_CP_676_elements(127) <= zeropad3D_CP_676_elements(126);
    -- CP-element group 128:  merge  place  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	499 
    -- CP-element group 128:  members (1) 
      -- CP-element group 128: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707__exit__
      -- 
    -- Element group zeropad3D_CP_676_elements(128) is bound as output of CP function.
    -- CP-element group 129:  merge  place  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	132 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_222/do_while_stmt_707/loop_back
      -- 
    -- Element group zeropad3D_CP_676_elements(129) is bound as output of CP function.
    -- CP-element group 130:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	135 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	497 
    -- CP-element group 130: 	498 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_222/do_while_stmt_707/condition_done
      -- CP-element group 130: 	 branch_block_stmt_222/do_while_stmt_707/loop_exit/$entry
      -- CP-element group 130: 	 branch_block_stmt_222/do_while_stmt_707/loop_taken/$entry
      -- 
    zeropad3D_CP_676_elements(130) <= zeropad3D_CP_676_elements(135);
    -- CP-element group 131:  branch  place  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	496 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (1) 
      -- CP-element group 131: 	 branch_block_stmt_222/do_while_stmt_707/loop_body_done
      -- 
    zeropad3D_CP_676_elements(131) <= zeropad3D_CP_676_elements(496);
    -- CP-element group 132:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	129 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	144 
    -- CP-element group 132: 	165 
    -- CP-element group 132: 	186 
    -- CP-element group 132:  members (1) 
      -- CP-element group 132: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/back_edge_to_loop_body
      -- 
    zeropad3D_CP_676_elements(132) <= zeropad3D_CP_676_elements(129);
    -- CP-element group 133:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	127 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	146 
    -- CP-element group 133: 	167 
    -- CP-element group 133: 	188 
    -- CP-element group 133:  members (1) 
      -- CP-element group 133: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/first_time_through_loop_body
      -- 
    zeropad3D_CP_676_elements(133) <= zeropad3D_CP_676_elements(127);
    -- CP-element group 134:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	140 
    -- CP-element group 134: 	141 
    -- CP-element group 134: 	159 
    -- CP-element group 134: 	160 
    -- CP-element group 134: 	333 
    -- CP-element group 134: 	369 
    -- CP-element group 134: 	180 
    -- CP-element group 134: 	181 
    -- CP-element group 134: 	410 
    -- CP-element group 134: 	411 
    -- CP-element group 134: 	441 
    -- CP-element group 134: 	442 
    -- CP-element group 134: 	476 
    -- CP-element group 134: 	477 
    -- CP-element group 134: 	494 
    -- CP-element group 134: 	205 
    -- CP-element group 134:  members (2) 
      -- CP-element group 134: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/loop_body_start
      -- CP-element group 134: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/$entry
      -- 
    -- Element group zeropad3D_CP_676_elements(134) is bound as output of CP function.
    -- CP-element group 135:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	139 
    -- CP-element group 135: 	316 
    -- CP-element group 135: 	494 
    -- CP-element group 135: 	256 
    -- CP-element group 135: 	264 
    -- CP-element group 135: 	268 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	130 
    -- CP-element group 135:  members (1) 
      -- CP-element group 135: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/condition_evaluated
      -- 
    condition_evaluated_1636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(135), ack => do_while_stmt_707_branch_req_0); -- 
    zeropad3D_cp_element_group_135: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_135"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(139) & zeropad3D_CP_676_elements(316) & zeropad3D_CP_676_elements(494) & zeropad3D_CP_676_elements(256) & zeropad3D_CP_676_elements(264) & zeropad3D_CP_676_elements(268);
      gj_zeropad3D_cp_element_group_135 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 136:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	140 
    -- CP-element group 136: 	159 
    -- CP-element group 136: 	180 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	139 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	161 
    -- CP-element group 136: 	182 
    -- CP-element group 136:  members (2) 
      -- CP-element group 136: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_709_sample_start__ps
      -- CP-element group 136: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/aggregated_phi_sample_req
      -- 
    zeropad3D_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(140) & zeropad3D_CP_676_elements(159) & zeropad3D_CP_676_elements(180) & zeropad3D_CP_676_elements(139);
      gj_zeropad3D_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	142 
    -- CP-element group 137: 	162 
    -- CP-element group 137: 	183 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	278 
    -- CP-element group 137: 	282 
    -- CP-element group 137: 	286 
    -- CP-element group 137: 	290 
    -- CP-element group 137: 	294 
    -- CP-element group 137: 	298 
    -- CP-element group 137: 	302 
    -- CP-element group 137: 	306 
    -- CP-element group 137: 	310 
    -- CP-element group 137: 	254 
    -- CP-element group 137: 	262 
    -- CP-element group 137: 	266 
    -- CP-element group 137: 	274 
    -- CP-element group 137: marked-successors 
    -- CP-element group 137: 	140 
    -- CP-element group 137: 	159 
    -- CP-element group 137: 	180 
    -- CP-element group 137:  members (4) 
      -- CP-element group 137: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_719_sample_completed_
      -- CP-element group 137: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_709_sample_completed_
      -- CP-element group 137: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_714_sample_completed_
      -- CP-element group 137: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/aggregated_phi_sample_ack
      -- 
    zeropad3D_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(142) & zeropad3D_CP_676_elements(162) & zeropad3D_CP_676_elements(183);
      gj_zeropad3D_cp_element_group_137 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	141 
    -- CP-element group 138: 	160 
    -- CP-element group 138: 	181 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	163 
    -- CP-element group 138: 	184 
    -- CP-element group 138:  members (2) 
      -- CP-element group 138: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_709_update_start__ps
      -- CP-element group 138: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/aggregated_phi_update_req
      -- 
    zeropad3D_cp_element_group_138: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_138"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(141) & zeropad3D_CP_676_elements(160) & zeropad3D_CP_676_elements(181);
      gj_zeropad3D_cp_element_group_138 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(138), clk => clk, reset => reset); --
    end block;
    -- CP-element group 139:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	143 
    -- CP-element group 139: 	164 
    -- CP-element group 139: 	185 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	135 
    -- CP-element group 139: marked-successors 
    -- CP-element group 139: 	136 
    -- CP-element group 139:  members (1) 
      -- CP-element group 139: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/aggregated_phi_update_ack
      -- 
    zeropad3D_cp_element_group_139: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_139"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(143) & zeropad3D_CP_676_elements(164) & zeropad3D_CP_676_elements(185);
      gj_zeropad3D_cp_element_group_139 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(139), clk => clk, reset => reset); --
    end block;
    -- CP-element group 140:  join  transition  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	134 
    -- CP-element group 140: marked-predecessors 
    -- CP-element group 140: 	276 
    -- CP-element group 140: 	280 
    -- CP-element group 140: 	137 
    -- CP-element group 140: 	256 
    -- CP-element group 140: 	264 
    -- CP-element group 140: 	268 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	136 
    -- CP-element group 140:  members (1) 
      -- CP-element group 140: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_709_sample_start_
      -- 
    zeropad3D_cp_element_group_140: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_140"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(134) & zeropad3D_CP_676_elements(276) & zeropad3D_CP_676_elements(280) & zeropad3D_CP_676_elements(137) & zeropad3D_CP_676_elements(256) & zeropad3D_CP_676_elements(264) & zeropad3D_CP_676_elements(268);
      gj_zeropad3D_cp_element_group_140 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(140), clk => clk, reset => reset); --
    end block;
    -- CP-element group 141:  join  transition  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	134 
    -- CP-element group 141: marked-predecessors 
    -- CP-element group 141: 	143 
    -- CP-element group 141: 	203 
    -- CP-element group 141: 	211 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	138 
    -- CP-element group 141:  members (1) 
      -- CP-element group 141: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_709_update_start_
      -- 
    zeropad3D_cp_element_group_141: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_141"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(134) & zeropad3D_CP_676_elements(143) & zeropad3D_CP_676_elements(203) & zeropad3D_CP_676_elements(211);
      gj_zeropad3D_cp_element_group_141 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(141), clk => clk, reset => reset); --
    end block;
    -- CP-element group 142:  join  transition  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	137 
    -- CP-element group 142:  members (1) 
      -- CP-element group 142: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_709_sample_completed__ps
      -- 
    -- Element group zeropad3D_CP_676_elements(142) is bound as output of CP function.
    -- CP-element group 143:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	139 
    -- CP-element group 143: 	201 
    -- CP-element group 143: 	209 
    -- CP-element group 143: marked-successors 
    -- CP-element group 143: 	141 
    -- CP-element group 143:  members (2) 
      -- CP-element group 143: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_709_update_completed__ps
      -- CP-element group 143: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_709_update_completed_
      -- 
    -- Element group zeropad3D_CP_676_elements(143) is bound as output of CP function.
    -- CP-element group 144:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	132 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (1) 
      -- CP-element group 144: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_709_loopback_trigger
      -- 
    zeropad3D_CP_676_elements(144) <= zeropad3D_CP_676_elements(132);
    -- CP-element group 145:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: successors 
    -- CP-element group 145:  members (2) 
      -- CP-element group 145: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_709_loopback_sample_req
      -- CP-element group 145: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_709_loopback_sample_req_ps
      -- 
    phi_stmt_709_loopback_sample_req_1651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_709_loopback_sample_req_1651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(145), ack => phi_stmt_709_req_0); -- 
    -- Element group zeropad3D_CP_676_elements(145) is bound as output of CP function.
    -- CP-element group 146:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	133 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (1) 
      -- CP-element group 146: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_709_entry_trigger
      -- 
    zeropad3D_CP_676_elements(146) <= zeropad3D_CP_676_elements(133);
    -- CP-element group 147:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (2) 
      -- CP-element group 147: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_709_entry_sample_req
      -- CP-element group 147: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_709_entry_sample_req_ps
      -- 
    phi_stmt_709_entry_sample_req_1654_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_709_entry_sample_req_1654_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(147), ack => phi_stmt_709_req_1); -- 
    -- Element group zeropad3D_CP_676_elements(147) is bound as output of CP function.
    -- CP-element group 148:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: successors 
    -- CP-element group 148:  members (2) 
      -- CP-element group 148: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_709_phi_mux_ack
      -- CP-element group 148: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_709_phi_mux_ack_ps
      -- 
    phi_stmt_709_phi_mux_ack_1657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_709_ack_0, ack => zeropad3D_CP_676_elements(148)); -- 
    -- CP-element group 149:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	151 
    -- CP-element group 149:  members (1) 
      -- CP-element group 149: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_712_sample_start__ps
      -- 
    -- Element group zeropad3D_CP_676_elements(149) is bound as output of CP function.
    -- CP-element group 150:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (1) 
      -- CP-element group 150: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_712_update_start__ps
      -- 
    -- Element group zeropad3D_CP_676_elements(150) is bound as output of CP function.
    -- CP-element group 151:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	149 
    -- CP-element group 151: marked-predecessors 
    -- CP-element group 151: 	153 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_712_sample_start_
      -- CP-element group 151: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_712_Sample/rr
      -- CP-element group 151: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_712_Sample/$entry
      -- 
    rr_1670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(151), ack => type_cast_712_inst_req_0); -- 
    zeropad3D_cp_element_group_151: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_151"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(149) & zeropad3D_CP_676_elements(153);
      gj_zeropad3D_cp_element_group_151 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(151), clk => clk, reset => reset); --
    end block;
    -- CP-element group 152:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: marked-predecessors 
    -- CP-element group 152: 	154 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	154 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_712_Update/cr
      -- CP-element group 152: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_712_Update/$entry
      -- CP-element group 152: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_712_update_start_
      -- 
    cr_1675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(152), ack => type_cast_712_inst_req_1); -- 
    zeropad3D_cp_element_group_152: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_152"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(150) & zeropad3D_CP_676_elements(154);
      gj_zeropad3D_cp_element_group_152 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(152), clk => clk, reset => reset); --
    end block;
    -- CP-element group 153:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153: marked-successors 
    -- CP-element group 153: 	151 
    -- CP-element group 153:  members (4) 
      -- CP-element group 153: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_712_Sample/$exit
      -- CP-element group 153: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_712_Sample/ra
      -- CP-element group 153: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_712_sample_completed__ps
      -- CP-element group 153: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_712_sample_completed_
      -- 
    ra_1671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_712_inst_ack_0, ack => zeropad3D_CP_676_elements(153)); -- 
    -- CP-element group 154:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	152 
    -- CP-element group 154: successors 
    -- CP-element group 154: marked-successors 
    -- CP-element group 154: 	152 
    -- CP-element group 154:  members (4) 
      -- CP-element group 154: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_712_Update/ca
      -- CP-element group 154: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_712_update_completed__ps
      -- CP-element group 154: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_712_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_712_Update/$exit
      -- 
    ca_1676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_712_inst_ack_1, ack => zeropad3D_CP_676_elements(154)); -- 
    -- CP-element group 155:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: successors 
    -- CP-element group 155:  members (4) 
      -- CP-element group 155: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/R_kx_x1_at_entry_713_sample_completed__ps
      -- CP-element group 155: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/R_kx_x1_at_entry_713_sample_start__ps
      -- CP-element group 155: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/R_kx_x1_at_entry_713_sample_completed_
      -- CP-element group 155: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/R_kx_x1_at_entry_713_sample_start_
      -- 
    -- Element group zeropad3D_CP_676_elements(155) is bound as output of CP function.
    -- CP-element group 156:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156:  members (2) 
      -- CP-element group 156: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/R_kx_x1_at_entry_713_update_start__ps
      -- CP-element group 156: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/R_kx_x1_at_entry_713_update_start_
      -- 
    -- Element group zeropad3D_CP_676_elements(156) is bound as output of CP function.
    -- CP-element group 157:  join  transition  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	158 
    -- CP-element group 157: successors 
    -- CP-element group 157:  members (1) 
      -- CP-element group 157: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/R_kx_x1_at_entry_713_update_completed__ps
      -- 
    zeropad3D_CP_676_elements(157) <= zeropad3D_CP_676_elements(158);
    -- CP-element group 158:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	156 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	157 
    -- CP-element group 158:  members (1) 
      -- CP-element group 158: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/R_kx_x1_at_entry_713_update_completed_
      -- 
    -- Element group zeropad3D_CP_676_elements(158) is a control-delay.
    cp_element_158_delay: control_delay_element  generic map(name => " 158_delay", delay_value => 1)  port map(req => zeropad3D_CP_676_elements(156), ack => zeropad3D_CP_676_elements(158), clk => clk, reset =>reset);
    -- CP-element group 159:  join  transition  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	134 
    -- CP-element group 159: marked-predecessors 
    -- CP-element group 159: 	137 
    -- CP-element group 159: 	284 
    -- CP-element group 159: 	288 
    -- CP-element group 159: 	292 
    -- CP-element group 159: 	296 
    -- CP-element group 159: 	256 
    -- CP-element group 159: 	264 
    -- CP-element group 159: 	268 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	136 
    -- CP-element group 159:  members (1) 
      -- CP-element group 159: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_714_sample_start_
      -- 
    zeropad3D_cp_element_group_159: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_159"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(134) & zeropad3D_CP_676_elements(137) & zeropad3D_CP_676_elements(284) & zeropad3D_CP_676_elements(288) & zeropad3D_CP_676_elements(292) & zeropad3D_CP_676_elements(296) & zeropad3D_CP_676_elements(256) & zeropad3D_CP_676_elements(264) & zeropad3D_CP_676_elements(268);
      gj_zeropad3D_cp_element_group_159 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(159), clk => clk, reset => reset); --
    end block;
    -- CP-element group 160:  join  transition  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	134 
    -- CP-element group 160: marked-predecessors 
    -- CP-element group 160: 	164 
    -- CP-element group 160: 	287 
    -- CP-element group 160: 	239 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	138 
    -- CP-element group 160:  members (1) 
      -- CP-element group 160: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_714_update_start_
      -- 
    zeropad3D_cp_element_group_160: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_160"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(134) & zeropad3D_CP_676_elements(164) & zeropad3D_CP_676_elements(287) & zeropad3D_CP_676_elements(239);
      gj_zeropad3D_cp_element_group_160 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(160), clk => clk, reset => reset); --
    end block;
    -- CP-element group 161:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	136 
    -- CP-element group 161: successors 
    -- CP-element group 161:  members (1) 
      -- CP-element group 161: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_714_sample_start__ps
      -- 
    zeropad3D_CP_676_elements(161) <= zeropad3D_CP_676_elements(136);
    -- CP-element group 162:  join  transition  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	137 
    -- CP-element group 162:  members (1) 
      -- CP-element group 162: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_714_sample_completed__ps
      -- 
    -- Element group zeropad3D_CP_676_elements(162) is bound as output of CP function.
    -- CP-element group 163:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	138 
    -- CP-element group 163: successors 
    -- CP-element group 163:  members (1) 
      -- CP-element group 163: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_714_update_start__ps
      -- 
    zeropad3D_CP_676_elements(163) <= zeropad3D_CP_676_elements(138);
    -- CP-element group 164:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	139 
    -- CP-element group 164: 	285 
    -- CP-element group 164: 	237 
    -- CP-element group 164: marked-successors 
    -- CP-element group 164: 	160 
    -- CP-element group 164:  members (2) 
      -- CP-element group 164: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_714_update_completed__ps
      -- CP-element group 164: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_714_update_completed_
      -- 
    -- Element group zeropad3D_CP_676_elements(164) is bound as output of CP function.
    -- CP-element group 165:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	132 
    -- CP-element group 165: successors 
    -- CP-element group 165:  members (1) 
      -- CP-element group 165: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_714_loopback_trigger
      -- 
    zeropad3D_CP_676_elements(165) <= zeropad3D_CP_676_elements(132);
    -- CP-element group 166:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: successors 
    -- CP-element group 166:  members (2) 
      -- CP-element group 166: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_714_loopback_sample_req
      -- CP-element group 166: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_714_loopback_sample_req_ps
      -- 
    phi_stmt_714_loopback_sample_req_1695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_714_loopback_sample_req_1695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(166), ack => phi_stmt_714_req_0); -- 
    -- Element group zeropad3D_CP_676_elements(166) is bound as output of CP function.
    -- CP-element group 167:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	133 
    -- CP-element group 167: successors 
    -- CP-element group 167:  members (1) 
      -- CP-element group 167: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_714_entry_trigger
      -- 
    zeropad3D_CP_676_elements(167) <= zeropad3D_CP_676_elements(133);
    -- CP-element group 168:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: successors 
    -- CP-element group 168:  members (2) 
      -- CP-element group 168: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_714_entry_sample_req_ps
      -- CP-element group 168: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_714_entry_sample_req
      -- 
    phi_stmt_714_entry_sample_req_1698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_714_entry_sample_req_1698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(168), ack => phi_stmt_714_req_1); -- 
    -- Element group zeropad3D_CP_676_elements(168) is bound as output of CP function.
    -- CP-element group 169:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: successors 
    -- CP-element group 169:  members (2) 
      -- CP-element group 169: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_714_phi_mux_ack_ps
      -- CP-element group 169: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_714_phi_mux_ack
      -- 
    phi_stmt_714_phi_mux_ack_1701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_714_ack_0, ack => zeropad3D_CP_676_elements(169)); -- 
    -- CP-element group 170:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	172 
    -- CP-element group 170:  members (1) 
      -- CP-element group 170: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_717_sample_start__ps
      -- 
    -- Element group zeropad3D_CP_676_elements(170) is bound as output of CP function.
    -- CP-element group 171:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	173 
    -- CP-element group 171:  members (1) 
      -- CP-element group 171: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_717_update_start__ps
      -- 
    -- Element group zeropad3D_CP_676_elements(171) is bound as output of CP function.
    -- CP-element group 172:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	170 
    -- CP-element group 172: marked-predecessors 
    -- CP-element group 172: 	174 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	174 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_717_Sample/rr
      -- CP-element group 172: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_717_Sample/$entry
      -- CP-element group 172: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_717_sample_start_
      -- 
    rr_1714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(172), ack => type_cast_717_inst_req_0); -- 
    zeropad3D_cp_element_group_172: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_172"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(170) & zeropad3D_CP_676_elements(174);
      gj_zeropad3D_cp_element_group_172 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(172), clk => clk, reset => reset); --
    end block;
    -- CP-element group 173:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	171 
    -- CP-element group 173: marked-predecessors 
    -- CP-element group 173: 	175 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	175 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_717_Update/cr
      -- CP-element group 173: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_717_Update/$entry
      -- CP-element group 173: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_717_update_start_
      -- 
    cr_1719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(173), ack => type_cast_717_inst_req_1); -- 
    zeropad3D_cp_element_group_173: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_173"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(171) & zeropad3D_CP_676_elements(175);
      gj_zeropad3D_cp_element_group_173 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(173), clk => clk, reset => reset); --
    end block;
    -- CP-element group 174:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	172 
    -- CP-element group 174: successors 
    -- CP-element group 174: marked-successors 
    -- CP-element group 174: 	172 
    -- CP-element group 174:  members (4) 
      -- CP-element group 174: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_717_Sample/ra
      -- CP-element group 174: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_717_Sample/$exit
      -- CP-element group 174: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_717_sample_completed_
      -- CP-element group 174: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_717_sample_completed__ps
      -- 
    ra_1715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_717_inst_ack_0, ack => zeropad3D_CP_676_elements(174)); -- 
    -- CP-element group 175:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	173 
    -- CP-element group 175: successors 
    -- CP-element group 175: marked-successors 
    -- CP-element group 175: 	173 
    -- CP-element group 175:  members (4) 
      -- CP-element group 175: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_717_Update/ca
      -- CP-element group 175: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_717_Update/$exit
      -- CP-element group 175: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_717_update_completed_
      -- CP-element group 175: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_717_update_completed__ps
      -- 
    ca_1720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_717_inst_ack_1, ack => zeropad3D_CP_676_elements(175)); -- 
    -- CP-element group 176:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: successors 
    -- CP-element group 176:  members (4) 
      -- CP-element group 176: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/R_i138x_x2_at_entry_718_sample_completed_
      -- CP-element group 176: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/R_i138x_x2_at_entry_718_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/R_i138x_x2_at_entry_718_sample_completed__ps
      -- CP-element group 176: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/R_i138x_x2_at_entry_718_sample_start__ps
      -- 
    -- Element group zeropad3D_CP_676_elements(176) is bound as output of CP function.
    -- CP-element group 177:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	179 
    -- CP-element group 177:  members (2) 
      -- CP-element group 177: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/R_i138x_x2_at_entry_718_update_start_
      -- CP-element group 177: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/R_i138x_x2_at_entry_718_update_start__ps
      -- 
    -- Element group zeropad3D_CP_676_elements(177) is bound as output of CP function.
    -- CP-element group 178:  join  transition  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	179 
    -- CP-element group 178: successors 
    -- CP-element group 178:  members (1) 
      -- CP-element group 178: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/R_i138x_x2_at_entry_718_update_completed__ps
      -- 
    zeropad3D_CP_676_elements(178) <= zeropad3D_CP_676_elements(179);
    -- CP-element group 179:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	177 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	178 
    -- CP-element group 179:  members (1) 
      -- CP-element group 179: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/R_i138x_x2_at_entry_718_update_completed_
      -- 
    -- Element group zeropad3D_CP_676_elements(179) is a control-delay.
    cp_element_179_delay: control_delay_element  generic map(name => " 179_delay", delay_value => 1)  port map(req => zeropad3D_CP_676_elements(177), ack => zeropad3D_CP_676_elements(179), clk => clk, reset =>reset);
    -- CP-element group 180:  join  transition  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	134 
    -- CP-element group 180: marked-predecessors 
    -- CP-element group 180: 	137 
    -- CP-element group 180: 	300 
    -- CP-element group 180: 	304 
    -- CP-element group 180: 	308 
    -- CP-element group 180: 	312 
    -- CP-element group 180: 	256 
    -- CP-element group 180: 	264 
    -- CP-element group 180: 	268 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	136 
    -- CP-element group 180:  members (1) 
      -- CP-element group 180: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_719_sample_start_
      -- 
    zeropad3D_cp_element_group_180: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_180"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(134) & zeropad3D_CP_676_elements(137) & zeropad3D_CP_676_elements(300) & zeropad3D_CP_676_elements(304) & zeropad3D_CP_676_elements(308) & zeropad3D_CP_676_elements(312) & zeropad3D_CP_676_elements(256) & zeropad3D_CP_676_elements(264) & zeropad3D_CP_676_elements(268);
      gj_zeropad3D_cp_element_group_180 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(180), clk => clk, reset => reset); --
    end block;
    -- CP-element group 181:  join  transition  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	134 
    -- CP-element group 181: marked-predecessors 
    -- CP-element group 181: 	185 
    -- CP-element group 181: 	303 
    -- CP-element group 181: 	215 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	138 
    -- CP-element group 181:  members (1) 
      -- CP-element group 181: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_719_update_start_
      -- 
    zeropad3D_cp_element_group_181: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_181"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(134) & zeropad3D_CP_676_elements(185) & zeropad3D_CP_676_elements(303) & zeropad3D_CP_676_elements(215);
      gj_zeropad3D_cp_element_group_181 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(181), clk => clk, reset => reset); --
    end block;
    -- CP-element group 182:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	136 
    -- CP-element group 182: successors 
    -- CP-element group 182:  members (1) 
      -- CP-element group 182: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_719_sample_start__ps
      -- 
    zeropad3D_CP_676_elements(182) <= zeropad3D_CP_676_elements(136);
    -- CP-element group 183:  join  transition  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	137 
    -- CP-element group 183:  members (1) 
      -- CP-element group 183: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_719_sample_completed__ps
      -- 
    -- Element group zeropad3D_CP_676_elements(183) is bound as output of CP function.
    -- CP-element group 184:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	138 
    -- CP-element group 184: successors 
    -- CP-element group 184:  members (1) 
      -- CP-element group 184: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_719_update_start__ps
      -- 
    zeropad3D_CP_676_elements(184) <= zeropad3D_CP_676_elements(138);
    -- CP-element group 185:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	139 
    -- CP-element group 185: 	301 
    -- CP-element group 185: 	213 
    -- CP-element group 185: marked-successors 
    -- CP-element group 185: 	181 
    -- CP-element group 185:  members (2) 
      -- CP-element group 185: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_719_update_completed_
      -- CP-element group 185: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_719_update_completed__ps
      -- 
    -- Element group zeropad3D_CP_676_elements(185) is bound as output of CP function.
    -- CP-element group 186:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	132 
    -- CP-element group 186: successors 
    -- CP-element group 186:  members (1) 
      -- CP-element group 186: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_719_loopback_trigger
      -- 
    zeropad3D_CP_676_elements(186) <= zeropad3D_CP_676_elements(132);
    -- CP-element group 187:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: successors 
    -- CP-element group 187:  members (2) 
      -- CP-element group 187: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_719_loopback_sample_req_ps
      -- CP-element group 187: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_719_loopback_sample_req
      -- 
    phi_stmt_719_loopback_sample_req_1739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_719_loopback_sample_req_1739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(187), ack => phi_stmt_719_req_0); -- 
    -- Element group zeropad3D_CP_676_elements(187) is bound as output of CP function.
    -- CP-element group 188:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	133 
    -- CP-element group 188: successors 
    -- CP-element group 188:  members (1) 
      -- CP-element group 188: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_719_entry_trigger
      -- 
    zeropad3D_CP_676_elements(188) <= zeropad3D_CP_676_elements(133);
    -- CP-element group 189:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: successors 
    -- CP-element group 189:  members (2) 
      -- CP-element group 189: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_719_entry_sample_req_ps
      -- CP-element group 189: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_719_entry_sample_req
      -- 
    phi_stmt_719_entry_sample_req_1742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_719_entry_sample_req_1742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(189), ack => phi_stmt_719_req_1); -- 
    -- Element group zeropad3D_CP_676_elements(189) is bound as output of CP function.
    -- CP-element group 190:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: successors 
    -- CP-element group 190:  members (2) 
      -- CP-element group 190: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_719_phi_mux_ack_ps
      -- CP-element group 190: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/phi_stmt_719_phi_mux_ack
      -- 
    phi_stmt_719_phi_mux_ack_1745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_719_ack_0, ack => zeropad3D_CP_676_elements(190)); -- 
    -- CP-element group 191:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	193 
    -- CP-element group 191:  members (1) 
      -- CP-element group 191: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_722_sample_start__ps
      -- 
    -- Element group zeropad3D_CP_676_elements(191) is bound as output of CP function.
    -- CP-element group 192:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	194 
    -- CP-element group 192:  members (1) 
      -- CP-element group 192: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_722_update_start__ps
      -- 
    -- Element group zeropad3D_CP_676_elements(192) is bound as output of CP function.
    -- CP-element group 193:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	191 
    -- CP-element group 193: marked-predecessors 
    -- CP-element group 193: 	195 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	195 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_722_sample_start_
      -- CP-element group 193: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_722_Sample/$entry
      -- CP-element group 193: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_722_Sample/rr
      -- 
    rr_1758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(193), ack => type_cast_722_inst_req_0); -- 
    zeropad3D_cp_element_group_193: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_193"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(191) & zeropad3D_CP_676_elements(195);
      gj_zeropad3D_cp_element_group_193 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(193), clk => clk, reset => reset); --
    end block;
    -- CP-element group 194:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	192 
    -- CP-element group 194: marked-predecessors 
    -- CP-element group 194: 	196 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	196 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_722_update_start_
      -- CP-element group 194: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_722_Update/$entry
      -- CP-element group 194: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_722_Update/cr
      -- 
    cr_1763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(194), ack => type_cast_722_inst_req_1); -- 
    zeropad3D_cp_element_group_194: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_194"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(192) & zeropad3D_CP_676_elements(196);
      gj_zeropad3D_cp_element_group_194 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(194), clk => clk, reset => reset); --
    end block;
    -- CP-element group 195:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	193 
    -- CP-element group 195: successors 
    -- CP-element group 195: marked-successors 
    -- CP-element group 195: 	193 
    -- CP-element group 195:  members (4) 
      -- CP-element group 195: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_722_sample_completed_
      -- CP-element group 195: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_722_sample_completed__ps
      -- CP-element group 195: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_722_Sample/$exit
      -- CP-element group 195: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_722_Sample/ra
      -- 
    ra_1759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_722_inst_ack_0, ack => zeropad3D_CP_676_elements(195)); -- 
    -- CP-element group 196:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	194 
    -- CP-element group 196: successors 
    -- CP-element group 196: marked-successors 
    -- CP-element group 196: 	194 
    -- CP-element group 196:  members (4) 
      -- CP-element group 196: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_722_update_completed__ps
      -- CP-element group 196: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_722_update_completed_
      -- CP-element group 196: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_722_Update/$exit
      -- CP-element group 196: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_722_Update/ca
      -- 
    ca_1764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_722_inst_ack_1, ack => zeropad3D_CP_676_elements(196)); -- 
    -- CP-element group 197:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: successors 
    -- CP-element group 197:  members (4) 
      -- CP-element group 197: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/R_jx_x1_at_entry_723_sample_completed_
      -- CP-element group 197: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/R_jx_x1_at_entry_723_sample_start_
      -- CP-element group 197: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/R_jx_x1_at_entry_723_sample_completed__ps
      -- CP-element group 197: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/R_jx_x1_at_entry_723_sample_start__ps
      -- 
    -- Element group zeropad3D_CP_676_elements(197) is bound as output of CP function.
    -- CP-element group 198:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	200 
    -- CP-element group 198:  members (2) 
      -- CP-element group 198: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/R_jx_x1_at_entry_723_update_start_
      -- CP-element group 198: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/R_jx_x1_at_entry_723_update_start__ps
      -- 
    -- Element group zeropad3D_CP_676_elements(198) is bound as output of CP function.
    -- CP-element group 199:  join  transition  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	200 
    -- CP-element group 199: successors 
    -- CP-element group 199:  members (1) 
      -- CP-element group 199: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/R_jx_x1_at_entry_723_update_completed__ps
      -- 
    zeropad3D_CP_676_elements(199) <= zeropad3D_CP_676_elements(200);
    -- CP-element group 200:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	198 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	199 
    -- CP-element group 200:  members (1) 
      -- CP-element group 200: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/R_jx_x1_at_entry_723_update_completed_
      -- 
    -- Element group zeropad3D_CP_676_elements(200) is a control-delay.
    cp_element_200_delay: control_delay_element  generic map(name => " 200_delay", delay_value => 1)  port map(req => zeropad3D_CP_676_elements(198), ack => zeropad3D_CP_676_elements(200), clk => clk, reset =>reset);
    -- CP-element group 201:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	143 
    -- CP-element group 201: marked-predecessors 
    -- CP-element group 201: 	203 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	203 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_727_Sample/rr
      -- CP-element group 201: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_727_Sample/$entry
      -- CP-element group 201: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_727_sample_start_
      -- 
    rr_1781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(201), ack => type_cast_727_inst_req_0); -- 
    zeropad3D_cp_element_group_201: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_201"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(143) & zeropad3D_CP_676_elements(203);
      gj_zeropad3D_cp_element_group_201 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(201), clk => clk, reset => reset); --
    end block;
    -- CP-element group 202:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: marked-predecessors 
    -- CP-element group 202: 	283 
    -- CP-element group 202: 	204 
    -- CP-element group 202: 	299 
    -- CP-element group 202: 	315 
    -- CP-element group 202: 	219 
    -- CP-element group 202: 	223 
    -- CP-element group 202: 	227 
    -- CP-element group 202: 	235 
    -- CP-element group 202: 	243 
    -- CP-element group 202: 	251 
    -- CP-element group 202: 	259 
    -- CP-element group 202: 	263 
    -- CP-element group 202: 	267 
    -- CP-element group 202: 	271 
    -- CP-element group 202: 	275 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	204 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_727_Update/cr
      -- CP-element group 202: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_727_Update/$entry
      -- CP-element group 202: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_727_update_start_
      -- 
    cr_1786_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1786_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(202), ack => type_cast_727_inst_req_1); -- 
    zeropad3D_cp_element_group_202: block -- 
      constant place_capacities: IntegerArray(0 to 14) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1);
      constant place_markings: IntegerArray(0 to 14)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1);
      constant place_delays: IntegerArray(0 to 14) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_202"; 
      signal preds: BooleanArray(1 to 15); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(283) & zeropad3D_CP_676_elements(204) & zeropad3D_CP_676_elements(299) & zeropad3D_CP_676_elements(315) & zeropad3D_CP_676_elements(219) & zeropad3D_CP_676_elements(223) & zeropad3D_CP_676_elements(227) & zeropad3D_CP_676_elements(235) & zeropad3D_CP_676_elements(243) & zeropad3D_CP_676_elements(251) & zeropad3D_CP_676_elements(259) & zeropad3D_CP_676_elements(263) & zeropad3D_CP_676_elements(267) & zeropad3D_CP_676_elements(271) & zeropad3D_CP_676_elements(275);
      gj_zeropad3D_cp_element_group_202 : generic_join generic map(name => joinName, number_of_predecessors => 15, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(202), clk => clk, reset => reset); --
    end block;
    -- CP-element group 203:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	201 
    -- CP-element group 203: successors 
    -- CP-element group 203: marked-successors 
    -- CP-element group 203: 	141 
    -- CP-element group 203: 	201 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_727_Sample/ra
      -- CP-element group 203: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_727_Sample/$exit
      -- CP-element group 203: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_727_sample_completed_
      -- 
    ra_1782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_727_inst_ack_0, ack => zeropad3D_CP_676_elements(203)); -- 
    -- CP-element group 204:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	202 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	281 
    -- CP-element group 204: 	297 
    -- CP-element group 204: 	313 
    -- CP-element group 204: 	217 
    -- CP-element group 204: 	221 
    -- CP-element group 204: 	225 
    -- CP-element group 204: 	233 
    -- CP-element group 204: 	241 
    -- CP-element group 204: 	249 
    -- CP-element group 204: 	257 
    -- CP-element group 204: 	261 
    -- CP-element group 204: 	265 
    -- CP-element group 204: 	269 
    -- CP-element group 204: 	273 
    -- CP-element group 204: marked-successors 
    -- CP-element group 204: 	202 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_727_Update/ca
      -- CP-element group 204: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_727_Update/$exit
      -- CP-element group 204: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_727_update_completed_
      -- 
    ca_1787_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_727_inst_ack_1, ack => zeropad3D_CP_676_elements(204)); -- 
    -- CP-element group 205:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	134 
    -- CP-element group 205: marked-predecessors 
    -- CP-element group 205: 	207 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	207 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_731_Sample/$entry
      -- CP-element group 205: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_731_sample_start_
      -- CP-element group 205: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_731_Sample/rr
      -- 
    rr_1795_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1795_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(205), ack => type_cast_731_inst_req_0); -- 
    zeropad3D_cp_element_group_205: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_205"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(134) & zeropad3D_CP_676_elements(207);
      gj_zeropad3D_cp_element_group_205 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(205), clk => clk, reset => reset); --
    end block;
    -- CP-element group 206:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: marked-predecessors 
    -- CP-element group 206: 	283 
    -- CP-element group 206: 	299 
    -- CP-element group 206: 	315 
    -- CP-element group 206: 	208 
    -- CP-element group 206: 	219 
    -- CP-element group 206: 	223 
    -- CP-element group 206: 	227 
    -- CP-element group 206: 	235 
    -- CP-element group 206: 	243 
    -- CP-element group 206: 	251 
    -- CP-element group 206: 	259 
    -- CP-element group 206: 	263 
    -- CP-element group 206: 	267 
    -- CP-element group 206: 	271 
    -- CP-element group 206: 	275 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	208 
    -- CP-element group 206:  members (3) 
      -- CP-element group 206: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_731_update_start_
      -- CP-element group 206: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_731_Update/cr
      -- CP-element group 206: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_731_Update/$entry
      -- 
    cr_1800_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1800_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(206), ack => type_cast_731_inst_req_1); -- 
    zeropad3D_cp_element_group_206: block -- 
      constant place_capacities: IntegerArray(0 to 14) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1);
      constant place_markings: IntegerArray(0 to 14)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1);
      constant place_delays: IntegerArray(0 to 14) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_206"; 
      signal preds: BooleanArray(1 to 15); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(283) & zeropad3D_CP_676_elements(299) & zeropad3D_CP_676_elements(315) & zeropad3D_CP_676_elements(208) & zeropad3D_CP_676_elements(219) & zeropad3D_CP_676_elements(223) & zeropad3D_CP_676_elements(227) & zeropad3D_CP_676_elements(235) & zeropad3D_CP_676_elements(243) & zeropad3D_CP_676_elements(251) & zeropad3D_CP_676_elements(259) & zeropad3D_CP_676_elements(263) & zeropad3D_CP_676_elements(267) & zeropad3D_CP_676_elements(271) & zeropad3D_CP_676_elements(275);
      gj_zeropad3D_cp_element_group_206 : generic_join generic map(name => joinName, number_of_predecessors => 15, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(206), clk => clk, reset => reset); --
    end block;
    -- CP-element group 207:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	205 
    -- CP-element group 207: successors 
    -- CP-element group 207: marked-successors 
    -- CP-element group 207: 	205 
    -- CP-element group 207:  members (3) 
      -- CP-element group 207: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_731_sample_completed_
      -- CP-element group 207: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_731_Sample/ra
      -- CP-element group 207: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_731_Sample/$exit
      -- 
    ra_1796_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_731_inst_ack_0, ack => zeropad3D_CP_676_elements(207)); -- 
    -- CP-element group 208:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	206 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	281 
    -- CP-element group 208: 	297 
    -- CP-element group 208: 	313 
    -- CP-element group 208: 	217 
    -- CP-element group 208: 	221 
    -- CP-element group 208: 	225 
    -- CP-element group 208: 	233 
    -- CP-element group 208: 	241 
    -- CP-element group 208: 	249 
    -- CP-element group 208: 	257 
    -- CP-element group 208: 	261 
    -- CP-element group 208: 	265 
    -- CP-element group 208: 	269 
    -- CP-element group 208: 	273 
    -- CP-element group 208: marked-successors 
    -- CP-element group 208: 	206 
    -- CP-element group 208:  members (3) 
      -- CP-element group 208: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_731_update_completed_
      -- CP-element group 208: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_731_Update/ca
      -- CP-element group 208: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_731_Update/$exit
      -- 
    ca_1801_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_731_inst_ack_1, ack => zeropad3D_CP_676_elements(208)); -- 
    -- CP-element group 209:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	143 
    -- CP-element group 209: marked-predecessors 
    -- CP-element group 209: 	211 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	211 
    -- CP-element group 209:  members (3) 
      -- CP-element group 209: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_751_Sample/$entry
      -- CP-element group 209: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_751_sample_start_
      -- CP-element group 209: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_751_Sample/req
      -- 
    req_1809_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1809_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(209), ack => W_kx_x1_748_delayed_1_0_749_inst_req_0); -- 
    zeropad3D_cp_element_group_209: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_209"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(143) & zeropad3D_CP_676_elements(211);
      gj_zeropad3D_cp_element_group_209 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(209), clk => clk, reset => reset); --
    end block;
    -- CP-element group 210:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: marked-predecessors 
    -- CP-element group 210: 	279 
    -- CP-element group 210: 	212 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	212 
    -- CP-element group 210:  members (3) 
      -- CP-element group 210: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_751_Update/req
      -- CP-element group 210: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_751_update_start_
      -- CP-element group 210: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_751_Update/$entry
      -- 
    req_1814_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1814_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(210), ack => W_kx_x1_748_delayed_1_0_749_inst_req_1); -- 
    zeropad3D_cp_element_group_210: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_210"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(279) & zeropad3D_CP_676_elements(212);
      gj_zeropad3D_cp_element_group_210 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(210), clk => clk, reset => reset); --
    end block;
    -- CP-element group 211:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	209 
    -- CP-element group 211: successors 
    -- CP-element group 211: marked-successors 
    -- CP-element group 211: 	141 
    -- CP-element group 211: 	209 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_751_Sample/$exit
      -- CP-element group 211: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_751_sample_completed_
      -- CP-element group 211: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_751_Sample/ack
      -- 
    ack_1810_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_kx_x1_748_delayed_1_0_749_inst_ack_0, ack => zeropad3D_CP_676_elements(211)); -- 
    -- CP-element group 212:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	210 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	277 
    -- CP-element group 212: marked-successors 
    -- CP-element group 212: 	210 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_751_Update/ack
      -- CP-element group 212: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_751_update_completed_
      -- CP-element group 212: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_751_Update/$exit
      -- 
    ack_1815_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_kx_x1_748_delayed_1_0_749_inst_ack_1, ack => zeropad3D_CP_676_elements(212)); -- 
    -- CP-element group 213:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	185 
    -- CP-element group 213: marked-predecessors 
    -- CP-element group 213: 	215 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	215 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_767_Sample/req
      -- CP-element group 213: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_767_Sample/$entry
      -- CP-element group 213: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_767_sample_start_
      -- 
    req_1823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(213), ack => W_jx_x1_761_delayed_1_0_765_inst_req_0); -- 
    zeropad3D_cp_element_group_213: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_213"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(185) & zeropad3D_CP_676_elements(215);
      gj_zeropad3D_cp_element_group_213 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(213), clk => clk, reset => reset); --
    end block;
    -- CP-element group 214:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: marked-predecessors 
    -- CP-element group 214: 	216 
    -- CP-element group 214: 	219 
    -- CP-element group 214: 	247 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	216 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_767_Update/req
      -- CP-element group 214: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_767_Update/$entry
      -- CP-element group 214: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_767_update_start_
      -- 
    req_1828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(214), ack => W_jx_x1_761_delayed_1_0_765_inst_req_1); -- 
    zeropad3D_cp_element_group_214: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_214"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(216) & zeropad3D_CP_676_elements(219) & zeropad3D_CP_676_elements(247);
      gj_zeropad3D_cp_element_group_214 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(214), clk => clk, reset => reset); --
    end block;
    -- CP-element group 215:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	213 
    -- CP-element group 215: successors 
    -- CP-element group 215: marked-successors 
    -- CP-element group 215: 	181 
    -- CP-element group 215: 	213 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_767_Sample/ack
      -- CP-element group 215: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_767_Sample/$exit
      -- CP-element group 215: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_767_sample_completed_
      -- 
    ack_1824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_jx_x1_761_delayed_1_0_765_inst_ack_0, ack => zeropad3D_CP_676_elements(215)); -- 
    -- CP-element group 216:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	214 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	217 
    -- CP-element group 216: 	245 
    -- CP-element group 216: marked-successors 
    -- CP-element group 216: 	214 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_767_Update/$exit
      -- CP-element group 216: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_767_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_767_Update/ack
      -- 
    ack_1829_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_jx_x1_761_delayed_1_0_765_inst_ack_1, ack => zeropad3D_CP_676_elements(216)); -- 
    -- CP-element group 217:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	204 
    -- CP-element group 217: 	208 
    -- CP-element group 217: 	216 
    -- CP-element group 217: marked-predecessors 
    -- CP-element group 217: 	219 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	219 
    -- CP-element group 217:  members (3) 
      -- CP-element group 217: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_778_sample_start_
      -- CP-element group 217: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_778_Sample/rr
      -- CP-element group 217: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_778_Sample/$entry
      -- 
    rr_1837_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1837_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(217), ack => type_cast_778_inst_req_0); -- 
    zeropad3D_cp_element_group_217: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_217"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(204) & zeropad3D_CP_676_elements(208) & zeropad3D_CP_676_elements(216) & zeropad3D_CP_676_elements(219);
      gj_zeropad3D_cp_element_group_217 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(217), clk => clk, reset => reset); --
    end block;
    -- CP-element group 218:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: marked-predecessors 
    -- CP-element group 218: 	307 
    -- CP-element group 218: 	311 
    -- CP-element group 218: 	220 
    -- CP-element group 218: 	231 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	220 
    -- CP-element group 218:  members (3) 
      -- CP-element group 218: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_778_update_start_
      -- CP-element group 218: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_778_Update/cr
      -- CP-element group 218: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_778_Update/$entry
      -- 
    cr_1842_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1842_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(218), ack => type_cast_778_inst_req_1); -- 
    zeropad3D_cp_element_group_218: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_218"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(307) & zeropad3D_CP_676_elements(311) & zeropad3D_CP_676_elements(220) & zeropad3D_CP_676_elements(231);
      gj_zeropad3D_cp_element_group_218 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(218), clk => clk, reset => reset); --
    end block;
    -- CP-element group 219:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	217 
    -- CP-element group 219: successors 
    -- CP-element group 219: marked-successors 
    -- CP-element group 219: 	202 
    -- CP-element group 219: 	206 
    -- CP-element group 219: 	214 
    -- CP-element group 219: 	217 
    -- CP-element group 219:  members (3) 
      -- CP-element group 219: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_778_sample_completed_
      -- CP-element group 219: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_778_Sample/ra
      -- CP-element group 219: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_778_Sample/$exit
      -- 
    ra_1838_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_778_inst_ack_0, ack => zeropad3D_CP_676_elements(219)); -- 
    -- CP-element group 220:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	218 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	305 
    -- CP-element group 220: 	309 
    -- CP-element group 220: 	229 
    -- CP-element group 220: marked-successors 
    -- CP-element group 220: 	218 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_778_update_completed_
      -- CP-element group 220: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_778_Update/ca
      -- CP-element group 220: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_778_Update/$exit
      -- 
    ca_1843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_778_inst_ack_1, ack => zeropad3D_CP_676_elements(220)); -- 
    -- CP-element group 221:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	204 
    -- CP-element group 221: 	208 
    -- CP-element group 221: marked-predecessors 
    -- CP-element group 221: 	223 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	223 
    -- CP-element group 221:  members (3) 
      -- CP-element group 221: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_782_sample_start_
      -- CP-element group 221: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_782_Sample/$entry
      -- CP-element group 221: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_782_Sample/req
      -- 
    req_1851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(221), ack => W_ifx_xelse_exec_guard_771_delayed_1_0_780_inst_req_0); -- 
    zeropad3D_cp_element_group_221: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_221"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(204) & zeropad3D_CP_676_elements(208) & zeropad3D_CP_676_elements(223);
      gj_zeropad3D_cp_element_group_221 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(221), clk => clk, reset => reset); --
    end block;
    -- CP-element group 222:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: marked-predecessors 
    -- CP-element group 222: 	224 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	224 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_782_update_start_
      -- CP-element group 222: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_782_Update/$entry
      -- CP-element group 222: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_782_Update/req
      -- 
    req_1856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(222), ack => W_ifx_xelse_exec_guard_771_delayed_1_0_780_inst_req_1); -- 
    zeropad3D_cp_element_group_222: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_222"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad3D_CP_676_elements(224);
      gj_zeropad3D_cp_element_group_222 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(222), clk => clk, reset => reset); --
    end block;
    -- CP-element group 223:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	221 
    -- CP-element group 223: successors 
    -- CP-element group 223: marked-successors 
    -- CP-element group 223: 	202 
    -- CP-element group 223: 	206 
    -- CP-element group 223: 	221 
    -- CP-element group 223:  members (3) 
      -- CP-element group 223: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_782_sample_completed_
      -- CP-element group 223: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_782_Sample/$exit
      -- CP-element group 223: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_782_Sample/ack
      -- 
    ack_1852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse_exec_guard_771_delayed_1_0_780_inst_ack_0, ack => zeropad3D_CP_676_elements(223)); -- 
    -- CP-element group 224:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	222 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	496 
    -- CP-element group 224: marked-successors 
    -- CP-element group 224: 	222 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_782_update_completed_
      -- CP-element group 224: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_782_Update/$exit
      -- CP-element group 224: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_782_Update/ack
      -- 
    ack_1857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse_exec_guard_771_delayed_1_0_780_inst_ack_1, ack => zeropad3D_CP_676_elements(224)); -- 
    -- CP-element group 225:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	204 
    -- CP-element group 225: 	208 
    -- CP-element group 225: marked-predecessors 
    -- CP-element group 225: 	227 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	227 
    -- CP-element group 225:  members (3) 
      -- CP-element group 225: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_791_sample_start_
      -- CP-element group 225: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_791_Sample/$entry
      -- CP-element group 225: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_791_Sample/req
      -- 
    req_1865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(225), ack => W_ifx_xelse_exec_guard_777_delayed_1_0_789_inst_req_0); -- 
    zeropad3D_cp_element_group_225: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_225"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(204) & zeropad3D_CP_676_elements(208) & zeropad3D_CP_676_elements(227);
      gj_zeropad3D_cp_element_group_225 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(225), clk => clk, reset => reset); --
    end block;
    -- CP-element group 226:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: marked-predecessors 
    -- CP-element group 226: 	228 
    -- CP-element group 226: 	231 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	228 
    -- CP-element group 226:  members (3) 
      -- CP-element group 226: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_791_update_start_
      -- CP-element group 226: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_791_Update/$entry
      -- CP-element group 226: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_791_Update/req
      -- 
    req_1870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(226), ack => W_ifx_xelse_exec_guard_777_delayed_1_0_789_inst_req_1); -- 
    zeropad3D_cp_element_group_226: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_226"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(228) & zeropad3D_CP_676_elements(231);
      gj_zeropad3D_cp_element_group_226 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(226), clk => clk, reset => reset); --
    end block;
    -- CP-element group 227:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	225 
    -- CP-element group 227: successors 
    -- CP-element group 227: marked-successors 
    -- CP-element group 227: 	202 
    -- CP-element group 227: 	206 
    -- CP-element group 227: 	225 
    -- CP-element group 227:  members (3) 
      -- CP-element group 227: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_791_sample_completed_
      -- CP-element group 227: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_791_Sample/$exit
      -- CP-element group 227: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_791_Sample/ack
      -- 
    ack_1866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse_exec_guard_777_delayed_1_0_789_inst_ack_0, ack => zeropad3D_CP_676_elements(227)); -- 
    -- CP-element group 228:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	226 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	229 
    -- CP-element group 228: marked-successors 
    -- CP-element group 228: 	226 
    -- CP-element group 228:  members (3) 
      -- CP-element group 228: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_791_update_completed_
      -- CP-element group 228: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_791_Update/$exit
      -- CP-element group 228: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_791_Update/ack
      -- 
    ack_1871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse_exec_guard_777_delayed_1_0_789_inst_ack_1, ack => zeropad3D_CP_676_elements(228)); -- 
    -- CP-element group 229:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	220 
    -- CP-element group 229: 	228 
    -- CP-element group 229: marked-predecessors 
    -- CP-element group 229: 	231 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	231 
    -- CP-element group 229:  members (3) 
      -- CP-element group 229: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_795_sample_start_
      -- CP-element group 229: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_795_Sample/$entry
      -- CP-element group 229: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_795_Sample/rr
      -- 
    rr_1879_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1879_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(229), ack => type_cast_795_inst_req_0); -- 
    zeropad3D_cp_element_group_229: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_229"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(220) & zeropad3D_CP_676_elements(228) & zeropad3D_CP_676_elements(231);
      gj_zeropad3D_cp_element_group_229 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(229), clk => clk, reset => reset); --
    end block;
    -- CP-element group 230:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: marked-predecessors 
    -- CP-element group 230: 	291 
    -- CP-element group 230: 	295 
    -- CP-element group 230: 	232 
    -- CP-element group 230: 	255 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	232 
    -- CP-element group 230:  members (3) 
      -- CP-element group 230: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_795_update_start_
      -- CP-element group 230: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_795_Update/$entry
      -- CP-element group 230: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_795_Update/cr
      -- 
    cr_1884_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1884_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(230), ack => type_cast_795_inst_req_1); -- 
    zeropad3D_cp_element_group_230: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_230"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(291) & zeropad3D_CP_676_elements(295) & zeropad3D_CP_676_elements(232) & zeropad3D_CP_676_elements(255);
      gj_zeropad3D_cp_element_group_230 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(230), clk => clk, reset => reset); --
    end block;
    -- CP-element group 231:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	229 
    -- CP-element group 231: successors 
    -- CP-element group 231: marked-successors 
    -- CP-element group 231: 	218 
    -- CP-element group 231: 	226 
    -- CP-element group 231: 	229 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_795_sample_completed_
      -- CP-element group 231: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_795_Sample/$exit
      -- CP-element group 231: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_795_Sample/ra
      -- 
    ra_1880_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_795_inst_ack_0, ack => zeropad3D_CP_676_elements(231)); -- 
    -- CP-element group 232:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	230 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	289 
    -- CP-element group 232: 	293 
    -- CP-element group 232: 	253 
    -- CP-element group 232: marked-successors 
    -- CP-element group 232: 	230 
    -- CP-element group 232:  members (3) 
      -- CP-element group 232: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_795_update_completed_
      -- CP-element group 232: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_795_Update/$exit
      -- CP-element group 232: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_795_Update/ca
      -- 
    ca_1885_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_795_inst_ack_1, ack => zeropad3D_CP_676_elements(232)); -- 
    -- CP-element group 233:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	204 
    -- CP-element group 233: 	208 
    -- CP-element group 233: marked-predecessors 
    -- CP-element group 233: 	235 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	235 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_799_sample_start_
      -- CP-element group 233: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_799_Sample/$entry
      -- CP-element group 233: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_799_Sample/req
      -- 
    req_1893_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1893_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(233), ack => W_ifx_xelse_exec_guard_782_delayed_2_0_797_inst_req_0); -- 
    zeropad3D_cp_element_group_233: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_233"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(204) & zeropad3D_CP_676_elements(208) & zeropad3D_CP_676_elements(235);
      gj_zeropad3D_cp_element_group_233 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(233), clk => clk, reset => reset); --
    end block;
    -- CP-element group 234:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: marked-predecessors 
    -- CP-element group 234: 	236 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	236 
    -- CP-element group 234:  members (3) 
      -- CP-element group 234: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_799_update_start_
      -- CP-element group 234: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_799_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_799_Update/req
      -- 
    req_1898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(234), ack => W_ifx_xelse_exec_guard_782_delayed_2_0_797_inst_req_1); -- 
    zeropad3D_cp_element_group_234: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_234"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad3D_CP_676_elements(236);
      gj_zeropad3D_cp_element_group_234 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(234), clk => clk, reset => reset); --
    end block;
    -- CP-element group 235:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	233 
    -- CP-element group 235: successors 
    -- CP-element group 235: marked-successors 
    -- CP-element group 235: 	202 
    -- CP-element group 235: 	206 
    -- CP-element group 235: 	233 
    -- CP-element group 235:  members (3) 
      -- CP-element group 235: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_799_sample_completed_
      -- CP-element group 235: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_799_Sample/$exit
      -- CP-element group 235: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_799_Sample/ack
      -- 
    ack_1894_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse_exec_guard_782_delayed_2_0_797_inst_ack_0, ack => zeropad3D_CP_676_elements(235)); -- 
    -- CP-element group 236:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	234 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	496 
    -- CP-element group 236: marked-successors 
    -- CP-element group 236: 	234 
    -- CP-element group 236:  members (3) 
      -- CP-element group 236: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_799_update_completed_
      -- CP-element group 236: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_799_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_799_Update/ack
      -- 
    ack_1899_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse_exec_guard_782_delayed_2_0_797_inst_ack_1, ack => zeropad3D_CP_676_elements(236)); -- 
    -- CP-element group 237:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	164 
    -- CP-element group 237: marked-predecessors 
    -- CP-element group 237: 	239 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	239 
    -- CP-element group 237:  members (3) 
      -- CP-element group 237: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_802_sample_start_
      -- CP-element group 237: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_802_Sample/$entry
      -- CP-element group 237: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_802_Sample/req
      -- 
    req_1907_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1907_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(237), ack => W_i138x_x2_785_delayed_3_0_800_inst_req_0); -- 
    zeropad3D_cp_element_group_237: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_237"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(164) & zeropad3D_CP_676_elements(239);
      gj_zeropad3D_cp_element_group_237 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(237), clk => clk, reset => reset); --
    end block;
    -- CP-element group 238:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: marked-predecessors 
    -- CP-element group 238: 	291 
    -- CP-element group 238: 	295 
    -- CP-element group 238: 	240 
    -- CP-element group 238: 	255 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	240 
    -- CP-element group 238:  members (3) 
      -- CP-element group 238: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_802_update_start_
      -- CP-element group 238: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_802_Update/$entry
      -- CP-element group 238: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_802_Update/req
      -- 
    req_1912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(238), ack => W_i138x_x2_785_delayed_3_0_800_inst_req_1); -- 
    zeropad3D_cp_element_group_238: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_238"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(291) & zeropad3D_CP_676_elements(295) & zeropad3D_CP_676_elements(240) & zeropad3D_CP_676_elements(255);
      gj_zeropad3D_cp_element_group_238 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(238), clk => clk, reset => reset); --
    end block;
    -- CP-element group 239:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	237 
    -- CP-element group 239: successors 
    -- CP-element group 239: marked-successors 
    -- CP-element group 239: 	160 
    -- CP-element group 239: 	237 
    -- CP-element group 239:  members (3) 
      -- CP-element group 239: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_802_sample_completed_
      -- CP-element group 239: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_802_Sample/$exit
      -- CP-element group 239: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_802_Sample/ack
      -- 
    ack_1908_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_i138x_x2_785_delayed_3_0_800_inst_ack_0, ack => zeropad3D_CP_676_elements(239)); -- 
    -- CP-element group 240:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	238 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	289 
    -- CP-element group 240: 	293 
    -- CP-element group 240: 	253 
    -- CP-element group 240: marked-successors 
    -- CP-element group 240: 	238 
    -- CP-element group 240:  members (3) 
      -- CP-element group 240: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_802_update_completed_
      -- CP-element group 240: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_802_Update/$exit
      -- CP-element group 240: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_802_Update/ack
      -- 
    ack_1913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_i138x_x2_785_delayed_3_0_800_inst_ack_1, ack => zeropad3D_CP_676_elements(240)); -- 
    -- CP-element group 241:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	204 
    -- CP-element group 241: 	208 
    -- CP-element group 241: marked-predecessors 
    -- CP-element group 241: 	243 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	243 
    -- CP-element group 241:  members (3) 
      -- CP-element group 241: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_811_sample_start_
      -- CP-element group 241: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_811_Sample/$entry
      -- CP-element group 241: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_811_Sample/req
      -- 
    req_1921_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1921_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(241), ack => W_ifx_xelse_exec_guard_788_delayed_1_0_809_inst_req_0); -- 
    zeropad3D_cp_element_group_241: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_241"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(204) & zeropad3D_CP_676_elements(208) & zeropad3D_CP_676_elements(243);
      gj_zeropad3D_cp_element_group_241 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(241), clk => clk, reset => reset); --
    end block;
    -- CP-element group 242:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: marked-predecessors 
    -- CP-element group 242: 	244 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	244 
    -- CP-element group 242:  members (3) 
      -- CP-element group 242: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_811_update_start_
      -- CP-element group 242: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_811_Update/$entry
      -- CP-element group 242: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_811_Update/req
      -- 
    req_1926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(242), ack => W_ifx_xelse_exec_guard_788_delayed_1_0_809_inst_req_1); -- 
    zeropad3D_cp_element_group_242: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_242"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad3D_CP_676_elements(244);
      gj_zeropad3D_cp_element_group_242 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(242), clk => clk, reset => reset); --
    end block;
    -- CP-element group 243:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	241 
    -- CP-element group 243: successors 
    -- CP-element group 243: marked-successors 
    -- CP-element group 243: 	202 
    -- CP-element group 243: 	206 
    -- CP-element group 243: 	241 
    -- CP-element group 243:  members (3) 
      -- CP-element group 243: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_811_sample_completed_
      -- CP-element group 243: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_811_Sample/$exit
      -- CP-element group 243: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_811_Sample/ack
      -- 
    ack_1922_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse_exec_guard_788_delayed_1_0_809_inst_ack_0, ack => zeropad3D_CP_676_elements(243)); -- 
    -- CP-element group 244:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	242 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	496 
    -- CP-element group 244: marked-successors 
    -- CP-element group 244: 	242 
    -- CP-element group 244:  members (3) 
      -- CP-element group 244: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_811_update_completed_
      -- CP-element group 244: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_811_Update/$exit
      -- CP-element group 244: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_811_Update/ack
      -- 
    ack_1927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse_exec_guard_788_delayed_1_0_809_inst_ack_1, ack => zeropad3D_CP_676_elements(244)); -- 
    -- CP-element group 245:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	216 
    -- CP-element group 245: marked-predecessors 
    -- CP-element group 245: 	247 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	247 
    -- CP-element group 245:  members (3) 
      -- CP-element group 245: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_814_sample_start_
      -- CP-element group 245: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_814_Sample/$entry
      -- CP-element group 245: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_814_Sample/req
      -- 
    req_1935_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1935_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(245), ack => W_inc187_793_delayed_1_0_812_inst_req_0); -- 
    zeropad3D_cp_element_group_245: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_245"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(216) & zeropad3D_CP_676_elements(247);
      gj_zeropad3D_cp_element_group_245 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(245), clk => clk, reset => reset); --
    end block;
    -- CP-element group 246:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: marked-predecessors 
    -- CP-element group 246: 	307 
    -- CP-element group 246: 	311 
    -- CP-element group 246: 	248 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	248 
    -- CP-element group 246:  members (3) 
      -- CP-element group 246: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_814_update_start_
      -- CP-element group 246: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_814_Update/$entry
      -- CP-element group 246: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_814_Update/req
      -- 
    req_1940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(246), ack => W_inc187_793_delayed_1_0_812_inst_req_1); -- 
    zeropad3D_cp_element_group_246: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_246"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(307) & zeropad3D_CP_676_elements(311) & zeropad3D_CP_676_elements(248);
      gj_zeropad3D_cp_element_group_246 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(246), clk => clk, reset => reset); --
    end block;
    -- CP-element group 247:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	245 
    -- CP-element group 247: successors 
    -- CP-element group 247: marked-successors 
    -- CP-element group 247: 	214 
    -- CP-element group 247: 	245 
    -- CP-element group 247:  members (3) 
      -- CP-element group 247: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_814_sample_completed_
      -- CP-element group 247: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_814_Sample/$exit
      -- CP-element group 247: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_814_Sample/ack
      -- 
    ack_1936_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_inc187_793_delayed_1_0_812_inst_ack_0, ack => zeropad3D_CP_676_elements(247)); -- 
    -- CP-element group 248:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	246 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	305 
    -- CP-element group 248: 	309 
    -- CP-element group 248: marked-successors 
    -- CP-element group 248: 	246 
    -- CP-element group 248:  members (3) 
      -- CP-element group 248: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_814_update_completed_
      -- CP-element group 248: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_814_Update/$exit
      -- CP-element group 248: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_814_Update/ack
      -- 
    ack_1941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_inc187_793_delayed_1_0_812_inst_ack_1, ack => zeropad3D_CP_676_elements(248)); -- 
    -- CP-element group 249:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	204 
    -- CP-element group 249: 	208 
    -- CP-element group 249: marked-predecessors 
    -- CP-element group 249: 	251 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	251 
    -- CP-element group 249:  members (3) 
      -- CP-element group 249: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_825_sample_start_
      -- CP-element group 249: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_825_Sample/$entry
      -- CP-element group 249: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_825_Sample/req
      -- 
    req_1949_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1949_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(249), ack => W_ifx_xelse_exec_guard_796_delayed_2_0_823_inst_req_0); -- 
    zeropad3D_cp_element_group_249: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_249"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(204) & zeropad3D_CP_676_elements(208) & zeropad3D_CP_676_elements(251);
      gj_zeropad3D_cp_element_group_249 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(249), clk => clk, reset => reset); --
    end block;
    -- CP-element group 250:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: marked-predecessors 
    -- CP-element group 250: 	252 
    -- CP-element group 250: 	255 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	252 
    -- CP-element group 250:  members (3) 
      -- CP-element group 250: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_825_update_start_
      -- CP-element group 250: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_825_Update/$entry
      -- CP-element group 250: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_825_Update/req
      -- 
    req_1954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(250), ack => W_ifx_xelse_exec_guard_796_delayed_2_0_823_inst_req_1); -- 
    zeropad3D_cp_element_group_250: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_250"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(252) & zeropad3D_CP_676_elements(255);
      gj_zeropad3D_cp_element_group_250 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(250), clk => clk, reset => reset); --
    end block;
    -- CP-element group 251:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	249 
    -- CP-element group 251: successors 
    -- CP-element group 251: marked-successors 
    -- CP-element group 251: 	202 
    -- CP-element group 251: 	206 
    -- CP-element group 251: 	249 
    -- CP-element group 251:  members (3) 
      -- CP-element group 251: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_825_sample_completed_
      -- CP-element group 251: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_825_Sample/$exit
      -- CP-element group 251: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_825_Sample/ack
      -- 
    ack_1950_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse_exec_guard_796_delayed_2_0_823_inst_ack_0, ack => zeropad3D_CP_676_elements(251)); -- 
    -- CP-element group 252:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	250 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	253 
    -- CP-element group 252: marked-successors 
    -- CP-element group 252: 	250 
    -- CP-element group 252:  members (3) 
      -- CP-element group 252: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_825_update_completed_
      -- CP-element group 252: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_825_Update/$exit
      -- CP-element group 252: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_825_Update/ack
      -- 
    ack_1955_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse_exec_guard_796_delayed_2_0_823_inst_ack_1, ack => zeropad3D_CP_676_elements(252)); -- 
    -- CP-element group 253:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	232 
    -- CP-element group 253: 	240 
    -- CP-element group 253: 	252 
    -- CP-element group 253: marked-predecessors 
    -- CP-element group 253: 	255 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	255 
    -- CP-element group 253:  members (3) 
      -- CP-element group 253: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_829_sample_start_
      -- CP-element group 253: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_829_Sample/$entry
      -- CP-element group 253: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_829_Sample/rr
      -- 
    rr_1963_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1963_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(253), ack => type_cast_829_inst_req_0); -- 
    zeropad3D_cp_element_group_253: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_253"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(232) & zeropad3D_CP_676_elements(240) & zeropad3D_CP_676_elements(252) & zeropad3D_CP_676_elements(255);
      gj_zeropad3D_cp_element_group_253 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(253), clk => clk, reset => reset); --
    end block;
    -- CP-element group 254:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	137 
    -- CP-element group 254: marked-predecessors 
    -- CP-element group 254: 	323 
    -- CP-element group 254: 	327 
    -- CP-element group 254: 	331 
    -- CP-element group 254: 	339 
    -- CP-element group 254: 	343 
    -- CP-element group 254: 	347 
    -- CP-element group 254: 	351 
    -- CP-element group 254: 	319 
    -- CP-element group 254: 	391 
    -- CP-element group 254: 	422 
    -- CP-element group 254: 	457 
    -- CP-element group 254: 	256 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	256 
    -- CP-element group 254:  members (3) 
      -- CP-element group 254: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_829_update_start_
      -- CP-element group 254: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_829_Update/$entry
      -- CP-element group 254: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_829_Update/cr
      -- 
    cr_1968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(254), ack => type_cast_829_inst_req_1); -- 
    zeropad3D_cp_element_group_254: block -- 
      constant place_capacities: IntegerArray(0 to 12) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1);
      constant place_markings: IntegerArray(0 to 12)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1);
      constant place_delays: IntegerArray(0 to 12) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_254"; 
      signal preds: BooleanArray(1 to 13); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(137) & zeropad3D_CP_676_elements(323) & zeropad3D_CP_676_elements(327) & zeropad3D_CP_676_elements(331) & zeropad3D_CP_676_elements(339) & zeropad3D_CP_676_elements(343) & zeropad3D_CP_676_elements(347) & zeropad3D_CP_676_elements(351) & zeropad3D_CP_676_elements(319) & zeropad3D_CP_676_elements(391) & zeropad3D_CP_676_elements(422) & zeropad3D_CP_676_elements(457) & zeropad3D_CP_676_elements(256);
      gj_zeropad3D_cp_element_group_254 : generic_join generic map(name => joinName, number_of_predecessors => 13, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(254), clk => clk, reset => reset); --
    end block;
    -- CP-element group 255:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	253 
    -- CP-element group 255: successors 
    -- CP-element group 255: marked-successors 
    -- CP-element group 255: 	230 
    -- CP-element group 255: 	238 
    -- CP-element group 255: 	250 
    -- CP-element group 255: 	253 
    -- CP-element group 255:  members (3) 
      -- CP-element group 255: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_829_sample_completed_
      -- CP-element group 255: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_829_Sample/$exit
      -- CP-element group 255: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_829_Sample/ra
      -- 
    ra_1964_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_829_inst_ack_0, ack => zeropad3D_CP_676_elements(255)); -- 
    -- CP-element group 256:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	254 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	135 
    -- CP-element group 256: 	325 
    -- CP-element group 256: 	329 
    -- CP-element group 256: 	337 
    -- CP-element group 256: 	341 
    -- CP-element group 256: 	345 
    -- CP-element group 256: 	349 
    -- CP-element group 256: 	317 
    -- CP-element group 256: 	321 
    -- CP-element group 256: 	389 
    -- CP-element group 256: 	420 
    -- CP-element group 256: 	455 
    -- CP-element group 256: marked-successors 
    -- CP-element group 256: 	140 
    -- CP-element group 256: 	159 
    -- CP-element group 256: 	180 
    -- CP-element group 256: 	254 
    -- CP-element group 256:  members (3) 
      -- CP-element group 256: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_829_update_completed_
      -- CP-element group 256: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_829_Update/$exit
      -- CP-element group 256: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_829_Update/ca
      -- 
    ca_1969_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_829_inst_ack_1, ack => zeropad3D_CP_676_elements(256)); -- 
    -- CP-element group 257:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	204 
    -- CP-element group 257: 	208 
    -- CP-element group 257: marked-predecessors 
    -- CP-element group 257: 	259 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	259 
    -- CP-element group 257:  members (3) 
      -- CP-element group 257: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_833_sample_start_
      -- CP-element group 257: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_833_Sample/$entry
      -- CP-element group 257: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_833_Sample/req
      -- 
    req_1977_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1977_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(257), ack => W_ifx_xelse_exec_guard_801_delayed_3_0_831_inst_req_0); -- 
    zeropad3D_cp_element_group_257: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_257"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(204) & zeropad3D_CP_676_elements(208) & zeropad3D_CP_676_elements(259);
      gj_zeropad3D_cp_element_group_257 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(257), clk => clk, reset => reset); --
    end block;
    -- CP-element group 258:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: marked-predecessors 
    -- CP-element group 258: 	260 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	260 
    -- CP-element group 258:  members (3) 
      -- CP-element group 258: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_833_update_start_
      -- CP-element group 258: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_833_Update/$entry
      -- CP-element group 258: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_833_Update/req
      -- 
    req_1982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(258), ack => W_ifx_xelse_exec_guard_801_delayed_3_0_831_inst_req_1); -- 
    zeropad3D_cp_element_group_258: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_258"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad3D_CP_676_elements(260);
      gj_zeropad3D_cp_element_group_258 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(258), clk => clk, reset => reset); --
    end block;
    -- CP-element group 259:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	257 
    -- CP-element group 259: successors 
    -- CP-element group 259: marked-successors 
    -- CP-element group 259: 	202 
    -- CP-element group 259: 	206 
    -- CP-element group 259: 	257 
    -- CP-element group 259:  members (3) 
      -- CP-element group 259: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_833_sample_completed_
      -- CP-element group 259: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_833_Sample/$exit
      -- CP-element group 259: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_833_Sample/ack
      -- 
    ack_1978_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse_exec_guard_801_delayed_3_0_831_inst_ack_0, ack => zeropad3D_CP_676_elements(259)); -- 
    -- CP-element group 260:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	258 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	496 
    -- CP-element group 260: marked-successors 
    -- CP-element group 260: 	258 
    -- CP-element group 260:  members (3) 
      -- CP-element group 260: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_833_update_completed_
      -- CP-element group 260: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_833_Update/$exit
      -- CP-element group 260: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_833_Update/ack
      -- 
    ack_1983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse_exec_guard_801_delayed_3_0_831_inst_ack_1, ack => zeropad3D_CP_676_elements(260)); -- 
    -- CP-element group 261:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	204 
    -- CP-element group 261: 	208 
    -- CP-element group 261: marked-predecessors 
    -- CP-element group 261: 	263 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	263 
    -- CP-element group 261:  members (3) 
      -- CP-element group 261: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_842_sample_start_
      -- CP-element group 261: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_842_Sample/$entry
      -- CP-element group 261: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_842_Sample/req
      -- 
    req_1991_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1991_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(261), ack => W_ifx_xelse_exec_guard_808_delayed_3_0_840_inst_req_0); -- 
    zeropad3D_cp_element_group_261: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_261"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(204) & zeropad3D_CP_676_elements(208) & zeropad3D_CP_676_elements(263);
      gj_zeropad3D_cp_element_group_261 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(261), clk => clk, reset => reset); --
    end block;
    -- CP-element group 262:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	137 
    -- CP-element group 262: marked-predecessors 
    -- CP-element group 262: 	323 
    -- CP-element group 262: 	327 
    -- CP-element group 262: 	331 
    -- CP-element group 262: 	339 
    -- CP-element group 262: 	343 
    -- CP-element group 262: 	347 
    -- CP-element group 262: 	351 
    -- CP-element group 262: 	319 
    -- CP-element group 262: 	391 
    -- CP-element group 262: 	422 
    -- CP-element group 262: 	457 
    -- CP-element group 262: 	264 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	264 
    -- CP-element group 262:  members (3) 
      -- CP-element group 262: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_842_update_start_
      -- CP-element group 262: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_842_Update/$entry
      -- CP-element group 262: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_842_Update/req
      -- 
    req_1996_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1996_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(262), ack => W_ifx_xelse_exec_guard_808_delayed_3_0_840_inst_req_1); -- 
    zeropad3D_cp_element_group_262: block -- 
      constant place_capacities: IntegerArray(0 to 12) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1);
      constant place_markings: IntegerArray(0 to 12)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1);
      constant place_delays: IntegerArray(0 to 12) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_262"; 
      signal preds: BooleanArray(1 to 13); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(137) & zeropad3D_CP_676_elements(323) & zeropad3D_CP_676_elements(327) & zeropad3D_CP_676_elements(331) & zeropad3D_CP_676_elements(339) & zeropad3D_CP_676_elements(343) & zeropad3D_CP_676_elements(347) & zeropad3D_CP_676_elements(351) & zeropad3D_CP_676_elements(319) & zeropad3D_CP_676_elements(391) & zeropad3D_CP_676_elements(422) & zeropad3D_CP_676_elements(457) & zeropad3D_CP_676_elements(264);
      gj_zeropad3D_cp_element_group_262 : generic_join generic map(name => joinName, number_of_predecessors => 13, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(262), clk => clk, reset => reset); --
    end block;
    -- CP-element group 263:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	261 
    -- CP-element group 263: successors 
    -- CP-element group 263: marked-successors 
    -- CP-element group 263: 	202 
    -- CP-element group 263: 	206 
    -- CP-element group 263: 	261 
    -- CP-element group 263:  members (3) 
      -- CP-element group 263: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_842_sample_completed_
      -- CP-element group 263: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_842_Sample/$exit
      -- CP-element group 263: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_842_Sample/ack
      -- 
    ack_1992_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse_exec_guard_808_delayed_3_0_840_inst_ack_0, ack => zeropad3D_CP_676_elements(263)); -- 
    -- CP-element group 264:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	262 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	135 
    -- CP-element group 264: 	325 
    -- CP-element group 264: 	329 
    -- CP-element group 264: 	337 
    -- CP-element group 264: 	341 
    -- CP-element group 264: 	345 
    -- CP-element group 264: 	349 
    -- CP-element group 264: 	317 
    -- CP-element group 264: 	321 
    -- CP-element group 264: 	389 
    -- CP-element group 264: 	420 
    -- CP-element group 264: 	455 
    -- CP-element group 264: marked-successors 
    -- CP-element group 264: 	140 
    -- CP-element group 264: 	159 
    -- CP-element group 264: 	180 
    -- CP-element group 264: 	262 
    -- CP-element group 264:  members (3) 
      -- CP-element group 264: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_842_update_completed_
      -- CP-element group 264: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_842_Update/$exit
      -- CP-element group 264: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_842_Update/ack
      -- 
    ack_1997_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse_exec_guard_808_delayed_3_0_840_inst_ack_1, ack => zeropad3D_CP_676_elements(264)); -- 
    -- CP-element group 265:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	204 
    -- CP-element group 265: 	208 
    -- CP-element group 265: marked-predecessors 
    -- CP-element group 265: 	267 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	267 
    -- CP-element group 265:  members (3) 
      -- CP-element group 265: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_850_sample_start_
      -- CP-element group 265: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_850_Sample/$entry
      -- CP-element group 265: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_850_Sample/req
      -- 
    req_2005_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2005_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(265), ack => W_ifx_xelse_exec_guard_813_delayed_3_0_848_inst_req_0); -- 
    zeropad3D_cp_element_group_265: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_265"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(204) & zeropad3D_CP_676_elements(208) & zeropad3D_CP_676_elements(267);
      gj_zeropad3D_cp_element_group_265 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(265), clk => clk, reset => reset); --
    end block;
    -- CP-element group 266:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	137 
    -- CP-element group 266: marked-predecessors 
    -- CP-element group 266: 	323 
    -- CP-element group 266: 	327 
    -- CP-element group 266: 	331 
    -- CP-element group 266: 	339 
    -- CP-element group 266: 	343 
    -- CP-element group 266: 	347 
    -- CP-element group 266: 	351 
    -- CP-element group 266: 	319 
    -- CP-element group 266: 	391 
    -- CP-element group 266: 	422 
    -- CP-element group 266: 	457 
    -- CP-element group 266: 	268 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	268 
    -- CP-element group 266:  members (3) 
      -- CP-element group 266: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_850_update_start_
      -- CP-element group 266: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_850_Update/$entry
      -- CP-element group 266: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_850_Update/req
      -- 
    req_2010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(266), ack => W_ifx_xelse_exec_guard_813_delayed_3_0_848_inst_req_1); -- 
    zeropad3D_cp_element_group_266: block -- 
      constant place_capacities: IntegerArray(0 to 12) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1);
      constant place_markings: IntegerArray(0 to 12)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1);
      constant place_delays: IntegerArray(0 to 12) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_266"; 
      signal preds: BooleanArray(1 to 13); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(137) & zeropad3D_CP_676_elements(323) & zeropad3D_CP_676_elements(327) & zeropad3D_CP_676_elements(331) & zeropad3D_CP_676_elements(339) & zeropad3D_CP_676_elements(343) & zeropad3D_CP_676_elements(347) & zeropad3D_CP_676_elements(351) & zeropad3D_CP_676_elements(319) & zeropad3D_CP_676_elements(391) & zeropad3D_CP_676_elements(422) & zeropad3D_CP_676_elements(457) & zeropad3D_CP_676_elements(268);
      gj_zeropad3D_cp_element_group_266 : generic_join generic map(name => joinName, number_of_predecessors => 13, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(266), clk => clk, reset => reset); --
    end block;
    -- CP-element group 267:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	265 
    -- CP-element group 267: successors 
    -- CP-element group 267: marked-successors 
    -- CP-element group 267: 	202 
    -- CP-element group 267: 	206 
    -- CP-element group 267: 	265 
    -- CP-element group 267:  members (3) 
      -- CP-element group 267: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_850_sample_completed_
      -- CP-element group 267: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_850_Sample/$exit
      -- CP-element group 267: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_850_Sample/ack
      -- 
    ack_2006_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse_exec_guard_813_delayed_3_0_848_inst_ack_0, ack => zeropad3D_CP_676_elements(267)); -- 
    -- CP-element group 268:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	266 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	135 
    -- CP-element group 268: 	325 
    -- CP-element group 268: 	329 
    -- CP-element group 268: 	337 
    -- CP-element group 268: 	341 
    -- CP-element group 268: 	345 
    -- CP-element group 268: 	349 
    -- CP-element group 268: 	317 
    -- CP-element group 268: 	321 
    -- CP-element group 268: 	389 
    -- CP-element group 268: 	420 
    -- CP-element group 268: 	455 
    -- CP-element group 268: marked-successors 
    -- CP-element group 268: 	140 
    -- CP-element group 268: 	159 
    -- CP-element group 268: 	180 
    -- CP-element group 268: 	266 
    -- CP-element group 268:  members (3) 
      -- CP-element group 268: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_850_update_completed_
      -- CP-element group 268: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_850_Update/$exit
      -- CP-element group 268: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_850_Update/ack
      -- 
    ack_2011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse_exec_guard_813_delayed_3_0_848_inst_ack_1, ack => zeropad3D_CP_676_elements(268)); -- 
    -- CP-element group 269:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	204 
    -- CP-element group 269: 	208 
    -- CP-element group 269: marked-predecessors 
    -- CP-element group 269: 	271 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	271 
    -- CP-element group 269:  members (3) 
      -- CP-element group 269: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_865_sample_start_
      -- CP-element group 269: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_865_Sample/$entry
      -- CP-element group 269: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_865_Sample/req
      -- 
    req_2019_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2019_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(269), ack => W_ifx_xthen_ifx_xend214_taken_826_delayed_3_0_863_inst_req_0); -- 
    zeropad3D_cp_element_group_269: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_269"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(204) & zeropad3D_CP_676_elements(208) & zeropad3D_CP_676_elements(271);
      gj_zeropad3D_cp_element_group_269 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(269), clk => clk, reset => reset); --
    end block;
    -- CP-element group 270:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: marked-predecessors 
    -- CP-element group 270: 	323 
    -- CP-element group 270: 	327 
    -- CP-element group 270: 	331 
    -- CP-element group 270: 	339 
    -- CP-element group 270: 	343 
    -- CP-element group 270: 	347 
    -- CP-element group 270: 	319 
    -- CP-element group 270: 	272 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	272 
    -- CP-element group 270:  members (3) 
      -- CP-element group 270: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_865_update_start_
      -- CP-element group 270: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_865_Update/$entry
      -- CP-element group 270: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_865_Update/req
      -- 
    req_2024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(270), ack => W_ifx_xthen_ifx_xend214_taken_826_delayed_3_0_863_inst_req_1); -- 
    zeropad3D_cp_element_group_270: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_270"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(323) & zeropad3D_CP_676_elements(327) & zeropad3D_CP_676_elements(331) & zeropad3D_CP_676_elements(339) & zeropad3D_CP_676_elements(343) & zeropad3D_CP_676_elements(347) & zeropad3D_CP_676_elements(319) & zeropad3D_CP_676_elements(272);
      gj_zeropad3D_cp_element_group_270 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(270), clk => clk, reset => reset); --
    end block;
    -- CP-element group 271:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	269 
    -- CP-element group 271: successors 
    -- CP-element group 271: marked-successors 
    -- CP-element group 271: 	202 
    -- CP-element group 271: 	206 
    -- CP-element group 271: 	269 
    -- CP-element group 271:  members (3) 
      -- CP-element group 271: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_865_sample_completed_
      -- CP-element group 271: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_865_Sample/$exit
      -- CP-element group 271: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_865_Sample/ack
      -- 
    ack_2020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen_ifx_xend214_taken_826_delayed_3_0_863_inst_ack_0, ack => zeropad3D_CP_676_elements(271)); -- 
    -- CP-element group 272:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	270 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	325 
    -- CP-element group 272: 	329 
    -- CP-element group 272: 	337 
    -- CP-element group 272: 	341 
    -- CP-element group 272: 	345 
    -- CP-element group 272: 	317 
    -- CP-element group 272: 	321 
    -- CP-element group 272: marked-successors 
    -- CP-element group 272: 	270 
    -- CP-element group 272:  members (3) 
      -- CP-element group 272: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_865_update_completed_
      -- CP-element group 272: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_865_Update/$exit
      -- CP-element group 272: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_865_Update/ack
      -- 
    ack_2025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen_ifx_xend214_taken_826_delayed_3_0_863_inst_ack_1, ack => zeropad3D_CP_676_elements(272)); -- 
    -- CP-element group 273:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	204 
    -- CP-element group 273: 	208 
    -- CP-element group 273: marked-predecessors 
    -- CP-element group 273: 	275 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	275 
    -- CP-element group 273:  members (3) 
      -- CP-element group 273: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_875_sample_start_
      -- CP-element group 273: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_875_Sample/$entry
      -- CP-element group 273: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_875_Sample/req
      -- 
    req_2033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(273), ack => W_ifx_xthen_ifx_xend214_taken_832_delayed_3_0_873_inst_req_0); -- 
    zeropad3D_cp_element_group_273: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_273"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(204) & zeropad3D_CP_676_elements(208) & zeropad3D_CP_676_elements(275);
      gj_zeropad3D_cp_element_group_273 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(273), clk => clk, reset => reset); --
    end block;
    -- CP-element group 274:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	137 
    -- CP-element group 274: marked-predecessors 
    -- CP-element group 274: 	276 
    -- CP-element group 274: 	391 
    -- CP-element group 274: 	422 
    -- CP-element group 274: 	457 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	276 
    -- CP-element group 274:  members (3) 
      -- CP-element group 274: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_875_update_start_
      -- CP-element group 274: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_875_Update/$entry
      -- CP-element group 274: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_875_Update/req
      -- 
    req_2038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(274), ack => W_ifx_xthen_ifx_xend214_taken_832_delayed_3_0_873_inst_req_1); -- 
    zeropad3D_cp_element_group_274: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_274"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(137) & zeropad3D_CP_676_elements(276) & zeropad3D_CP_676_elements(391) & zeropad3D_CP_676_elements(422) & zeropad3D_CP_676_elements(457);
      gj_zeropad3D_cp_element_group_274 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(274), clk => clk, reset => reset); --
    end block;
    -- CP-element group 275:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	273 
    -- CP-element group 275: successors 
    -- CP-element group 275: marked-successors 
    -- CP-element group 275: 	202 
    -- CP-element group 275: 	206 
    -- CP-element group 275: 	273 
    -- CP-element group 275:  members (3) 
      -- CP-element group 275: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_875_sample_completed_
      -- CP-element group 275: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_875_Sample/$exit
      -- CP-element group 275: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_875_Sample/ack
      -- 
    ack_2034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen_ifx_xend214_taken_832_delayed_3_0_873_inst_ack_0, ack => zeropad3D_CP_676_elements(275)); -- 
    -- CP-element group 276:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	274 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	389 
    -- CP-element group 276: 	420 
    -- CP-element group 276: 	455 
    -- CP-element group 276: marked-successors 
    -- CP-element group 276: 	140 
    -- CP-element group 276: 	274 
    -- CP-element group 276:  members (3) 
      -- CP-element group 276: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_875_update_completed_
      -- CP-element group 276: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_875_Update/$exit
      -- CP-element group 276: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_875_Update/ack
      -- 
    ack_2039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen_ifx_xend214_taken_832_delayed_3_0_873_inst_ack_1, ack => zeropad3D_CP_676_elements(276)); -- 
    -- CP-element group 277:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	212 
    -- CP-element group 277: marked-predecessors 
    -- CP-element group 277: 	279 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	279 
    -- CP-element group 277:  members (3) 
      -- CP-element group 277: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_878_sample_start_
      -- CP-element group 277: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_878_Sample/$entry
      -- CP-element group 277: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_878_Sample/rr
      -- 
    rr_2047_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2047_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(277), ack => type_cast_878_inst_req_0); -- 
    zeropad3D_cp_element_group_277: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_277"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(212) & zeropad3D_CP_676_elements(279);
      gj_zeropad3D_cp_element_group_277 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(277), clk => clk, reset => reset); --
    end block;
    -- CP-element group 278:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	137 
    -- CP-element group 278: marked-predecessors 
    -- CP-element group 278: 	280 
    -- CP-element group 278: 	391 
    -- CP-element group 278: 	422 
    -- CP-element group 278: 	457 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	280 
    -- CP-element group 278:  members (3) 
      -- CP-element group 278: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_878_update_start_
      -- CP-element group 278: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_878_Update/$entry
      -- CP-element group 278: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_878_Update/cr
      -- 
    cr_2052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(278), ack => type_cast_878_inst_req_1); -- 
    zeropad3D_cp_element_group_278: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_278"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(137) & zeropad3D_CP_676_elements(280) & zeropad3D_CP_676_elements(391) & zeropad3D_CP_676_elements(422) & zeropad3D_CP_676_elements(457);
      gj_zeropad3D_cp_element_group_278 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(278), clk => clk, reset => reset); --
    end block;
    -- CP-element group 279:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	277 
    -- CP-element group 279: successors 
    -- CP-element group 279: marked-successors 
    -- CP-element group 279: 	277 
    -- CP-element group 279: 	210 
    -- CP-element group 279:  members (3) 
      -- CP-element group 279: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_878_sample_completed_
      -- CP-element group 279: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_878_Sample/$exit
      -- CP-element group 279: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_878_Sample/ra
      -- 
    ra_2048_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_878_inst_ack_0, ack => zeropad3D_CP_676_elements(279)); -- 
    -- CP-element group 280:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	278 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	389 
    -- CP-element group 280: 	420 
    -- CP-element group 280: 	455 
    -- CP-element group 280: marked-successors 
    -- CP-element group 280: 	278 
    -- CP-element group 280: 	140 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_878_update_completed_
      -- CP-element group 280: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_878_Update/$exit
      -- CP-element group 280: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_878_Update/ca
      -- 
    ca_2053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_878_inst_ack_1, ack => zeropad3D_CP_676_elements(280)); -- 
    -- CP-element group 281:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	204 
    -- CP-element group 281: 	208 
    -- CP-element group 281: marked-predecessors 
    -- CP-element group 281: 	283 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	283 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_899_sample_start_
      -- CP-element group 281: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_899_Sample/$entry
      -- CP-element group 281: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_899_Sample/req
      -- 
    req_2061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(281), ack => W_ifx_xthen_ifx_xend214_taken_850_delayed_3_0_897_inst_req_0); -- 
    zeropad3D_cp_element_group_281: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_281"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(204) & zeropad3D_CP_676_elements(208) & zeropad3D_CP_676_elements(283);
      gj_zeropad3D_cp_element_group_281 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(281), clk => clk, reset => reset); --
    end block;
    -- CP-element group 282:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	137 
    -- CP-element group 282: marked-predecessors 
    -- CP-element group 282: 	319 
    -- CP-element group 282: 	391 
    -- CP-element group 282: 	284 
    -- CP-element group 282: 	422 
    -- CP-element group 282: 	457 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	284 
    -- CP-element group 282:  members (3) 
      -- CP-element group 282: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_899_update_start_
      -- CP-element group 282: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_899_Update/$entry
      -- CP-element group 282: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_899_Update/req
      -- 
    req_2066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(282), ack => W_ifx_xthen_ifx_xend214_taken_850_delayed_3_0_897_inst_req_1); -- 
    zeropad3D_cp_element_group_282: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_282"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(137) & zeropad3D_CP_676_elements(319) & zeropad3D_CP_676_elements(391) & zeropad3D_CP_676_elements(284) & zeropad3D_CP_676_elements(422) & zeropad3D_CP_676_elements(457);
      gj_zeropad3D_cp_element_group_282 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(282), clk => clk, reset => reset); --
    end block;
    -- CP-element group 283:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	281 
    -- CP-element group 283: successors 
    -- CP-element group 283: marked-successors 
    -- CP-element group 283: 	281 
    -- CP-element group 283: 	202 
    -- CP-element group 283: 	206 
    -- CP-element group 283:  members (3) 
      -- CP-element group 283: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_899_sample_completed_
      -- CP-element group 283: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_899_Sample/$exit
      -- CP-element group 283: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_899_Sample/ack
      -- 
    ack_2062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 283_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen_ifx_xend214_taken_850_delayed_3_0_897_inst_ack_0, ack => zeropad3D_CP_676_elements(283)); -- 
    -- CP-element group 284:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	282 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	317 
    -- CP-element group 284: 	389 
    -- CP-element group 284: 	420 
    -- CP-element group 284: 	455 
    -- CP-element group 284: marked-successors 
    -- CP-element group 284: 	282 
    -- CP-element group 284: 	159 
    -- CP-element group 284:  members (3) 
      -- CP-element group 284: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_899_update_completed_
      -- CP-element group 284: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_899_Update/$exit
      -- CP-element group 284: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_899_Update/ack
      -- 
    ack_2067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen_ifx_xend214_taken_850_delayed_3_0_897_inst_ack_1, ack => zeropad3D_CP_676_elements(284)); -- 
    -- CP-element group 285:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	164 
    -- CP-element group 285: marked-predecessors 
    -- CP-element group 285: 	287 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	287 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_902_sample_start_
      -- CP-element group 285: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_902_Sample/$entry
      -- CP-element group 285: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_902_Sample/rr
      -- 
    rr_2075_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2075_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(285), ack => type_cast_902_inst_req_0); -- 
    zeropad3D_cp_element_group_285: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_285"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(164) & zeropad3D_CP_676_elements(287);
      gj_zeropad3D_cp_element_group_285 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(285), clk => clk, reset => reset); --
    end block;
    -- CP-element group 286:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	137 
    -- CP-element group 286: marked-predecessors 
    -- CP-element group 286: 	319 
    -- CP-element group 286: 	391 
    -- CP-element group 286: 	422 
    -- CP-element group 286: 	288 
    -- CP-element group 286: 	457 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	288 
    -- CP-element group 286:  members (3) 
      -- CP-element group 286: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_902_update_start_
      -- CP-element group 286: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_902_Update/$entry
      -- CP-element group 286: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_902_Update/cr
      -- 
    cr_2080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(286), ack => type_cast_902_inst_req_1); -- 
    zeropad3D_cp_element_group_286: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_286"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(137) & zeropad3D_CP_676_elements(319) & zeropad3D_CP_676_elements(391) & zeropad3D_CP_676_elements(422) & zeropad3D_CP_676_elements(288) & zeropad3D_CP_676_elements(457);
      gj_zeropad3D_cp_element_group_286 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(286), clk => clk, reset => reset); --
    end block;
    -- CP-element group 287:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	285 
    -- CP-element group 287: successors 
    -- CP-element group 287: marked-successors 
    -- CP-element group 287: 	160 
    -- CP-element group 287: 	285 
    -- CP-element group 287:  members (3) 
      -- CP-element group 287: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_902_sample_completed_
      -- CP-element group 287: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_902_Sample/$exit
      -- CP-element group 287: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_902_Sample/ra
      -- 
    ra_2076_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_902_inst_ack_0, ack => zeropad3D_CP_676_elements(287)); -- 
    -- CP-element group 288:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	286 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	317 
    -- CP-element group 288: 	389 
    -- CP-element group 288: 	420 
    -- CP-element group 288: 	455 
    -- CP-element group 288: marked-successors 
    -- CP-element group 288: 	159 
    -- CP-element group 288: 	286 
    -- CP-element group 288:  members (3) 
      -- CP-element group 288: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_902_update_completed_
      -- CP-element group 288: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_902_Update/$exit
      -- CP-element group 288: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_902_Update/ca
      -- 
    ca_2081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_902_inst_ack_1, ack => zeropad3D_CP_676_elements(288)); -- 
    -- CP-element group 289:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	232 
    -- CP-element group 289: 	240 
    -- CP-element group 289: marked-predecessors 
    -- CP-element group 289: 	291 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	291 
    -- CP-element group 289:  members (3) 
      -- CP-element group 289: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_906_sample_start_
      -- CP-element group 289: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_906_Sample/$entry
      -- CP-element group 289: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_906_Sample/rr
      -- 
    rr_2089_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2089_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(289), ack => type_cast_906_inst_req_0); -- 
    zeropad3D_cp_element_group_289: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_289"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(232) & zeropad3D_CP_676_elements(240) & zeropad3D_CP_676_elements(291);
      gj_zeropad3D_cp_element_group_289 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(289), clk => clk, reset => reset); --
    end block;
    -- CP-element group 290:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	137 
    -- CP-element group 290: marked-predecessors 
    -- CP-element group 290: 	319 
    -- CP-element group 290: 	391 
    -- CP-element group 290: 	422 
    -- CP-element group 290: 	292 
    -- CP-element group 290: 	457 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	292 
    -- CP-element group 290:  members (3) 
      -- CP-element group 290: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_906_update_start_
      -- CP-element group 290: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_906_Update/$entry
      -- CP-element group 290: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_906_Update/cr
      -- 
    cr_2094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(290), ack => type_cast_906_inst_req_1); -- 
    zeropad3D_cp_element_group_290: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_290"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(137) & zeropad3D_CP_676_elements(319) & zeropad3D_CP_676_elements(391) & zeropad3D_CP_676_elements(422) & zeropad3D_CP_676_elements(292) & zeropad3D_CP_676_elements(457);
      gj_zeropad3D_cp_element_group_290 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(290), clk => clk, reset => reset); --
    end block;
    -- CP-element group 291:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	289 
    -- CP-element group 291: successors 
    -- CP-element group 291: marked-successors 
    -- CP-element group 291: 	289 
    -- CP-element group 291: 	230 
    -- CP-element group 291: 	238 
    -- CP-element group 291:  members (3) 
      -- CP-element group 291: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_906_sample_completed_
      -- CP-element group 291: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_906_Sample/$exit
      -- CP-element group 291: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_906_Sample/ra
      -- 
    ra_2090_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_906_inst_ack_0, ack => zeropad3D_CP_676_elements(291)); -- 
    -- CP-element group 292:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	290 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	317 
    -- CP-element group 292: 	389 
    -- CP-element group 292: 	420 
    -- CP-element group 292: 	455 
    -- CP-element group 292: marked-successors 
    -- CP-element group 292: 	159 
    -- CP-element group 292: 	290 
    -- CP-element group 292:  members (3) 
      -- CP-element group 292: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_906_update_completed_
      -- CP-element group 292: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_906_Update/$exit
      -- CP-element group 292: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_906_Update/ca
      -- 
    ca_2095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_906_inst_ack_1, ack => zeropad3D_CP_676_elements(292)); -- 
    -- CP-element group 293:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	232 
    -- CP-element group 293: 	240 
    -- CP-element group 293: marked-predecessors 
    -- CP-element group 293: 	295 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	295 
    -- CP-element group 293:  members (3) 
      -- CP-element group 293: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_910_sample_start_
      -- CP-element group 293: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_910_Sample/$entry
      -- CP-element group 293: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_910_Sample/rr
      -- 
    rr_2103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(293), ack => type_cast_910_inst_req_0); -- 
    zeropad3D_cp_element_group_293: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_293"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(232) & zeropad3D_CP_676_elements(240) & zeropad3D_CP_676_elements(295);
      gj_zeropad3D_cp_element_group_293 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(293), clk => clk, reset => reset); --
    end block;
    -- CP-element group 294:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	137 
    -- CP-element group 294: marked-predecessors 
    -- CP-element group 294: 	319 
    -- CP-element group 294: 	391 
    -- CP-element group 294: 	422 
    -- CP-element group 294: 	457 
    -- CP-element group 294: 	296 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	296 
    -- CP-element group 294:  members (3) 
      -- CP-element group 294: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_910_update_start_
      -- CP-element group 294: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_910_Update/$entry
      -- CP-element group 294: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_910_Update/cr
      -- 
    cr_2108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(294), ack => type_cast_910_inst_req_1); -- 
    zeropad3D_cp_element_group_294: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_294"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(137) & zeropad3D_CP_676_elements(319) & zeropad3D_CP_676_elements(391) & zeropad3D_CP_676_elements(422) & zeropad3D_CP_676_elements(457) & zeropad3D_CP_676_elements(296);
      gj_zeropad3D_cp_element_group_294 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(294), clk => clk, reset => reset); --
    end block;
    -- CP-element group 295:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	293 
    -- CP-element group 295: successors 
    -- CP-element group 295: marked-successors 
    -- CP-element group 295: 	293 
    -- CP-element group 295: 	230 
    -- CP-element group 295: 	238 
    -- CP-element group 295:  members (3) 
      -- CP-element group 295: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_910_sample_completed_
      -- CP-element group 295: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_910_Sample/$exit
      -- CP-element group 295: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_910_Sample/ra
      -- 
    ra_2104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_910_inst_ack_0, ack => zeropad3D_CP_676_elements(295)); -- 
    -- CP-element group 296:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	294 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	317 
    -- CP-element group 296: 	389 
    -- CP-element group 296: 	420 
    -- CP-element group 296: 	455 
    -- CP-element group 296: marked-successors 
    -- CP-element group 296: 	159 
    -- CP-element group 296: 	294 
    -- CP-element group 296:  members (3) 
      -- CP-element group 296: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_910_update_completed_
      -- CP-element group 296: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_910_Update/$exit
      -- CP-element group 296: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_910_Update/ca
      -- 
    ca_2109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_910_inst_ack_1, ack => zeropad3D_CP_676_elements(296)); -- 
    -- CP-element group 297:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	204 
    -- CP-element group 297: 	208 
    -- CP-element group 297: marked-predecessors 
    -- CP-element group 297: 	299 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	299 
    -- CP-element group 297:  members (3) 
      -- CP-element group 297: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_927_Sample/$entry
      -- CP-element group 297: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_927_Sample/req
      -- CP-element group 297: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_927_sample_start_
      -- 
    req_2117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(297), ack => W_ifx_xthen_ifx_xend214_taken_866_delayed_3_0_925_inst_req_0); -- 
    zeropad3D_cp_element_group_297: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_297"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(204) & zeropad3D_CP_676_elements(208) & zeropad3D_CP_676_elements(299);
      gj_zeropad3D_cp_element_group_297 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(297), clk => clk, reset => reset); --
    end block;
    -- CP-element group 298:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	137 
    -- CP-element group 298: marked-predecessors 
    -- CP-element group 298: 	351 
    -- CP-element group 298: 	391 
    -- CP-element group 298: 	422 
    -- CP-element group 298: 	457 
    -- CP-element group 298: 	300 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	300 
    -- CP-element group 298:  members (3) 
      -- CP-element group 298: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_927_Update/$entry
      -- CP-element group 298: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_927_update_start_
      -- CP-element group 298: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_927_Update/req
      -- 
    req_2122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(298), ack => W_ifx_xthen_ifx_xend214_taken_866_delayed_3_0_925_inst_req_1); -- 
    zeropad3D_cp_element_group_298: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_298"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(137) & zeropad3D_CP_676_elements(351) & zeropad3D_CP_676_elements(391) & zeropad3D_CP_676_elements(422) & zeropad3D_CP_676_elements(457) & zeropad3D_CP_676_elements(300);
      gj_zeropad3D_cp_element_group_298 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(298), clk => clk, reset => reset); --
    end block;
    -- CP-element group 299:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	297 
    -- CP-element group 299: successors 
    -- CP-element group 299: marked-successors 
    -- CP-element group 299: 	202 
    -- CP-element group 299: 	297 
    -- CP-element group 299: 	206 
    -- CP-element group 299:  members (3) 
      -- CP-element group 299: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_927_Sample/$exit
      -- CP-element group 299: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_927_Sample/ack
      -- CP-element group 299: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_927_sample_completed_
      -- 
    ack_2118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen_ifx_xend214_taken_866_delayed_3_0_925_inst_ack_0, ack => zeropad3D_CP_676_elements(299)); -- 
    -- CP-element group 300:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	298 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	349 
    -- CP-element group 300: 	389 
    -- CP-element group 300: 	420 
    -- CP-element group 300: 	455 
    -- CP-element group 300: marked-successors 
    -- CP-element group 300: 	180 
    -- CP-element group 300: 	298 
    -- CP-element group 300:  members (3) 
      -- CP-element group 300: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_927_Update/ack
      -- CP-element group 300: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_927_Update/$exit
      -- CP-element group 300: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_927_update_completed_
      -- 
    ack_2123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen_ifx_xend214_taken_866_delayed_3_0_925_inst_ack_1, ack => zeropad3D_CP_676_elements(300)); -- 
    -- CP-element group 301:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	185 
    -- CP-element group 301: marked-predecessors 
    -- CP-element group 301: 	303 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	303 
    -- CP-element group 301:  members (3) 
      -- CP-element group 301: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_930_sample_start_
      -- CP-element group 301: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_930_Sample/$entry
      -- CP-element group 301: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_930_Sample/rr
      -- 
    rr_2131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(301), ack => type_cast_930_inst_req_0); -- 
    zeropad3D_cp_element_group_301: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_301"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(185) & zeropad3D_CP_676_elements(303);
      gj_zeropad3D_cp_element_group_301 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(301), clk => clk, reset => reset); --
    end block;
    -- CP-element group 302:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	137 
    -- CP-element group 302: marked-predecessors 
    -- CP-element group 302: 	351 
    -- CP-element group 302: 	391 
    -- CP-element group 302: 	422 
    -- CP-element group 302: 	457 
    -- CP-element group 302: 	304 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	304 
    -- CP-element group 302:  members (3) 
      -- CP-element group 302: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_930_Update/$entry
      -- CP-element group 302: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_930_update_start_
      -- CP-element group 302: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_930_Update/cr
      -- 
    cr_2136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(302), ack => type_cast_930_inst_req_1); -- 
    zeropad3D_cp_element_group_302: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_302"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(137) & zeropad3D_CP_676_elements(351) & zeropad3D_CP_676_elements(391) & zeropad3D_CP_676_elements(422) & zeropad3D_CP_676_elements(457) & zeropad3D_CP_676_elements(304);
      gj_zeropad3D_cp_element_group_302 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(302), clk => clk, reset => reset); --
    end block;
    -- CP-element group 303:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	301 
    -- CP-element group 303: successors 
    -- CP-element group 303: marked-successors 
    -- CP-element group 303: 	181 
    -- CP-element group 303: 	301 
    -- CP-element group 303:  members (3) 
      -- CP-element group 303: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_930_sample_completed_
      -- CP-element group 303: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_930_Sample/$exit
      -- CP-element group 303: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_930_Sample/ra
      -- 
    ra_2132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_930_inst_ack_0, ack => zeropad3D_CP_676_elements(303)); -- 
    -- CP-element group 304:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	302 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	349 
    -- CP-element group 304: 	389 
    -- CP-element group 304: 	420 
    -- CP-element group 304: 	455 
    -- CP-element group 304: marked-successors 
    -- CP-element group 304: 	180 
    -- CP-element group 304: 	302 
    -- CP-element group 304:  members (3) 
      -- CP-element group 304: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_930_Update/ca
      -- CP-element group 304: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_930_Update/$exit
      -- CP-element group 304: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_930_update_completed_
      -- 
    ca_2137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_930_inst_ack_1, ack => zeropad3D_CP_676_elements(304)); -- 
    -- CP-element group 305:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	220 
    -- CP-element group 305: 	248 
    -- CP-element group 305: marked-predecessors 
    -- CP-element group 305: 	307 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	307 
    -- CP-element group 305:  members (3) 
      -- CP-element group 305: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_934_Sample/rr
      -- CP-element group 305: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_934_sample_start_
      -- CP-element group 305: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_934_Sample/$entry
      -- 
    rr_2145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(305), ack => type_cast_934_inst_req_0); -- 
    zeropad3D_cp_element_group_305: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_305"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(220) & zeropad3D_CP_676_elements(248) & zeropad3D_CP_676_elements(307);
      gj_zeropad3D_cp_element_group_305 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(305), clk => clk, reset => reset); --
    end block;
    -- CP-element group 306:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	137 
    -- CP-element group 306: marked-predecessors 
    -- CP-element group 306: 	351 
    -- CP-element group 306: 	391 
    -- CP-element group 306: 	422 
    -- CP-element group 306: 	457 
    -- CP-element group 306: 	308 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	308 
    -- CP-element group 306:  members (3) 
      -- CP-element group 306: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_934_update_start_
      -- CP-element group 306: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_934_Update/cr
      -- CP-element group 306: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_934_Update/$entry
      -- 
    cr_2150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(306), ack => type_cast_934_inst_req_1); -- 
    zeropad3D_cp_element_group_306: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_306"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(137) & zeropad3D_CP_676_elements(351) & zeropad3D_CP_676_elements(391) & zeropad3D_CP_676_elements(422) & zeropad3D_CP_676_elements(457) & zeropad3D_CP_676_elements(308);
      gj_zeropad3D_cp_element_group_306 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(306), clk => clk, reset => reset); --
    end block;
    -- CP-element group 307:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	305 
    -- CP-element group 307: successors 
    -- CP-element group 307: marked-successors 
    -- CP-element group 307: 	305 
    -- CP-element group 307: 	218 
    -- CP-element group 307: 	246 
    -- CP-element group 307:  members (3) 
      -- CP-element group 307: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_934_sample_completed_
      -- CP-element group 307: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_934_Sample/$exit
      -- CP-element group 307: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_934_Sample/ra
      -- 
    ra_2146_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_934_inst_ack_0, ack => zeropad3D_CP_676_elements(307)); -- 
    -- CP-element group 308:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	306 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	349 
    -- CP-element group 308: 	389 
    -- CP-element group 308: 	420 
    -- CP-element group 308: 	455 
    -- CP-element group 308: marked-successors 
    -- CP-element group 308: 	180 
    -- CP-element group 308: 	306 
    -- CP-element group 308:  members (3) 
      -- CP-element group 308: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_934_Update/ca
      -- CP-element group 308: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_934_update_completed_
      -- CP-element group 308: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_934_Update/$exit
      -- 
    ca_2151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_934_inst_ack_1, ack => zeropad3D_CP_676_elements(308)); -- 
    -- CP-element group 309:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	220 
    -- CP-element group 309: 	248 
    -- CP-element group 309: marked-predecessors 
    -- CP-element group 309: 	311 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	311 
    -- CP-element group 309:  members (3) 
      -- CP-element group 309: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_938_Sample/rr
      -- CP-element group 309: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_938_Sample/$entry
      -- CP-element group 309: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_938_sample_start_
      -- 
    rr_2159_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2159_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(309), ack => type_cast_938_inst_req_0); -- 
    zeropad3D_cp_element_group_309: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_309"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(220) & zeropad3D_CP_676_elements(248) & zeropad3D_CP_676_elements(311);
      gj_zeropad3D_cp_element_group_309 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(309), clk => clk, reset => reset); --
    end block;
    -- CP-element group 310:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	137 
    -- CP-element group 310: marked-predecessors 
    -- CP-element group 310: 	351 
    -- CP-element group 310: 	391 
    -- CP-element group 310: 	422 
    -- CP-element group 310: 	457 
    -- CP-element group 310: 	312 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	312 
    -- CP-element group 310:  members (3) 
      -- CP-element group 310: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_938_update_start_
      -- CP-element group 310: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_938_Update/$entry
      -- CP-element group 310: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_938_Update/cr
      -- 
    cr_2164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(310), ack => type_cast_938_inst_req_1); -- 
    zeropad3D_cp_element_group_310: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_310"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(137) & zeropad3D_CP_676_elements(351) & zeropad3D_CP_676_elements(391) & zeropad3D_CP_676_elements(422) & zeropad3D_CP_676_elements(457) & zeropad3D_CP_676_elements(312);
      gj_zeropad3D_cp_element_group_310 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(310), clk => clk, reset => reset); --
    end block;
    -- CP-element group 311:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	309 
    -- CP-element group 311: successors 
    -- CP-element group 311: marked-successors 
    -- CP-element group 311: 	309 
    -- CP-element group 311: 	218 
    -- CP-element group 311: 	246 
    -- CP-element group 311:  members (3) 
      -- CP-element group 311: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_938_Sample/$exit
      -- CP-element group 311: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_938_Sample/ra
      -- CP-element group 311: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_938_sample_completed_
      -- 
    ra_2160_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_938_inst_ack_0, ack => zeropad3D_CP_676_elements(311)); -- 
    -- CP-element group 312:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	310 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	349 
    -- CP-element group 312: 	389 
    -- CP-element group 312: 	420 
    -- CP-element group 312: 	455 
    -- CP-element group 312: marked-successors 
    -- CP-element group 312: 	180 
    -- CP-element group 312: 	310 
    -- CP-element group 312:  members (3) 
      -- CP-element group 312: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_938_update_completed_
      -- CP-element group 312: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_938_Update/$exit
      -- CP-element group 312: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_938_Update/ca
      -- 
    ca_2165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_938_inst_ack_1, ack => zeropad3D_CP_676_elements(312)); -- 
    -- CP-element group 313:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	204 
    -- CP-element group 313: 	208 
    -- CP-element group 313: marked-predecessors 
    -- CP-element group 313: 	315 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	315 
    -- CP-element group 313:  members (3) 
      -- CP-element group 313: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_955_sample_start_
      -- CP-element group 313: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_955_Sample/$entry
      -- CP-element group 313: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_955_Sample/req
      -- 
    req_2173_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2173_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(313), ack => W_ifx_xthen_ifx_xend214_taken_882_delayed_3_0_953_inst_req_0); -- 
    zeropad3D_cp_element_group_313: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_313"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(204) & zeropad3D_CP_676_elements(208) & zeropad3D_CP_676_elements(315);
      gj_zeropad3D_cp_element_group_313 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(313), clk => clk, reset => reset); --
    end block;
    -- CP-element group 314:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: marked-predecessors 
    -- CP-element group 314: 	316 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	316 
    -- CP-element group 314:  members (3) 
      -- CP-element group 314: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_955_update_start_
      -- CP-element group 314: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_955_Update/req
      -- CP-element group 314: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_955_Update/$entry
      -- 
    req_2178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(314), ack => W_ifx_xthen_ifx_xend214_taken_882_delayed_3_0_953_inst_req_1); -- 
    zeropad3D_cp_element_group_314: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_314"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad3D_CP_676_elements(316);
      gj_zeropad3D_cp_element_group_314 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(314), clk => clk, reset => reset); --
    end block;
    -- CP-element group 315:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	313 
    -- CP-element group 315: successors 
    -- CP-element group 315: marked-successors 
    -- CP-element group 315: 	202 
    -- CP-element group 315: 	206 
    -- CP-element group 315: 	313 
    -- CP-element group 315:  members (3) 
      -- CP-element group 315: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_955_sample_completed_
      -- CP-element group 315: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_955_Sample/$exit
      -- CP-element group 315: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_955_Sample/ack
      -- 
    ack_2174_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen_ifx_xend214_taken_882_delayed_3_0_953_inst_ack_0, ack => zeropad3D_CP_676_elements(315)); -- 
    -- CP-element group 316:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	314 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	135 
    -- CP-element group 316: marked-successors 
    -- CP-element group 316: 	314 
    -- CP-element group 316:  members (3) 
      -- CP-element group 316: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_955_Update/ack
      -- CP-element group 316: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_955_update_completed_
      -- CP-element group 316: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_955_Update/$exit
      -- 
    ack_2179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen_ifx_xend214_taken_882_delayed_3_0_953_inst_ack_1, ack => zeropad3D_CP_676_elements(316)); -- 
    -- CP-element group 317:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	284 
    -- CP-element group 317: 	288 
    -- CP-element group 317: 	292 
    -- CP-element group 317: 	296 
    -- CP-element group 317: 	256 
    -- CP-element group 317: 	264 
    -- CP-element group 317: 	268 
    -- CP-element group 317: 	272 
    -- CP-element group 317: marked-predecessors 
    -- CP-element group 317: 	319 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	319 
    -- CP-element group 317:  members (3) 
      -- CP-element group 317: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1038_Sample/$entry
      -- CP-element group 317: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1038_Sample/rr
      -- CP-element group 317: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1038_sample_start_
      -- 
    rr_2187_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2187_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(317), ack => type_cast_1038_inst_req_0); -- 
    zeropad3D_cp_element_group_317: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 1);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_317"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(284) & zeropad3D_CP_676_elements(288) & zeropad3D_CP_676_elements(292) & zeropad3D_CP_676_elements(296) & zeropad3D_CP_676_elements(256) & zeropad3D_CP_676_elements(264) & zeropad3D_CP_676_elements(268) & zeropad3D_CP_676_elements(272) & zeropad3D_CP_676_elements(319);
      gj_zeropad3D_cp_element_group_317 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(317), clk => clk, reset => reset); --
    end block;
    -- CP-element group 318:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: marked-predecessors 
    -- CP-element group 318: 	355 
    -- CP-element group 318: 	359 
    -- CP-element group 318: 	363 
    -- CP-element group 318: 	320 
    -- CP-element group 318: 	367 
    -- CP-element group 318: 	375 
    -- CP-element group 318: 	379 
    -- CP-element group 318: 	383 
    -- CP-element group 318: 	387 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	320 
    -- CP-element group 318:  members (3) 
      -- CP-element group 318: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1038_update_start_
      -- CP-element group 318: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1038_Update/cr
      -- CP-element group 318: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1038_Update/$entry
      -- 
    cr_2192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(318), ack => type_cast_1038_inst_req_1); -- 
    zeropad3D_cp_element_group_318: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_318"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(355) & zeropad3D_CP_676_elements(359) & zeropad3D_CP_676_elements(363) & zeropad3D_CP_676_elements(320) & zeropad3D_CP_676_elements(367) & zeropad3D_CP_676_elements(375) & zeropad3D_CP_676_elements(379) & zeropad3D_CP_676_elements(383) & zeropad3D_CP_676_elements(387);
      gj_zeropad3D_cp_element_group_318 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(318), clk => clk, reset => reset); --
    end block;
    -- CP-element group 319:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	317 
    -- CP-element group 319: successors 
    -- CP-element group 319: marked-successors 
    -- CP-element group 319: 	282 
    -- CP-element group 319: 	317 
    -- CP-element group 319: 	286 
    -- CP-element group 319: 	290 
    -- CP-element group 319: 	294 
    -- CP-element group 319: 	254 
    -- CP-element group 319: 	262 
    -- CP-element group 319: 	266 
    -- CP-element group 319: 	270 
    -- CP-element group 319:  members (3) 
      -- CP-element group 319: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1038_sample_completed_
      -- CP-element group 319: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1038_Sample/$exit
      -- CP-element group 319: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1038_Sample/ra
      -- 
    ra_2188_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 319_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1038_inst_ack_0, ack => zeropad3D_CP_676_elements(319)); -- 
    -- CP-element group 320:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	318 
    -- CP-element group 320: successors 
    -- CP-element group 320: 	353 
    -- CP-element group 320: 	357 
    -- CP-element group 320: 	361 
    -- CP-element group 320: 	365 
    -- CP-element group 320: 	373 
    -- CP-element group 320: 	377 
    -- CP-element group 320: 	381 
    -- CP-element group 320: 	385 
    -- CP-element group 320: marked-successors 
    -- CP-element group 320: 	318 
    -- CP-element group 320:  members (3) 
      -- CP-element group 320: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1038_Update/ca
      -- CP-element group 320: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1038_update_completed_
      -- CP-element group 320: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1038_Update/$exit
      -- 
    ca_2193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 320_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1038_inst_ack_1, ack => zeropad3D_CP_676_elements(320)); -- 
    -- CP-element group 321:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	256 
    -- CP-element group 321: 	264 
    -- CP-element group 321: 	268 
    -- CP-element group 321: 	272 
    -- CP-element group 321: marked-predecessors 
    -- CP-element group 321: 	323 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	323 
    -- CP-element group 321:  members (3) 
      -- CP-element group 321: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1042_sample_start_
      -- CP-element group 321: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1042_Sample/req
      -- CP-element group 321: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1042_Sample/$entry
      -- 
    req_2201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(321), ack => W_ifx_xend214_exec_guard_965_delayed_1_0_1040_inst_req_0); -- 
    zeropad3D_cp_element_group_321: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_321"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(256) & zeropad3D_CP_676_elements(264) & zeropad3D_CP_676_elements(268) & zeropad3D_CP_676_elements(272) & zeropad3D_CP_676_elements(323);
      gj_zeropad3D_cp_element_group_321 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(321), clk => clk, reset => reset); --
    end block;
    -- CP-element group 322:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: marked-predecessors 
    -- CP-element group 322: 	324 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	324 
    -- CP-element group 322:  members (3) 
      -- CP-element group 322: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1042_update_start_
      -- CP-element group 322: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1042_Update/req
      -- CP-element group 322: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1042_Update/$entry
      -- 
    req_2206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(322), ack => W_ifx_xend214_exec_guard_965_delayed_1_0_1040_inst_req_1); -- 
    zeropad3D_cp_element_group_322: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_322"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad3D_CP_676_elements(324);
      gj_zeropad3D_cp_element_group_322 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(322), clk => clk, reset => reset); --
    end block;
    -- CP-element group 323:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	321 
    -- CP-element group 323: successors 
    -- CP-element group 323: marked-successors 
    -- CP-element group 323: 	321 
    -- CP-element group 323: 	254 
    -- CP-element group 323: 	262 
    -- CP-element group 323: 	266 
    -- CP-element group 323: 	270 
    -- CP-element group 323:  members (3) 
      -- CP-element group 323: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1042_sample_completed_
      -- CP-element group 323: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1042_Sample/ack
      -- CP-element group 323: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1042_Sample/$exit
      -- 
    ack_2202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 323_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend214_exec_guard_965_delayed_1_0_1040_inst_ack_0, ack => zeropad3D_CP_676_elements(323)); -- 
    -- CP-element group 324:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	322 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	496 
    -- CP-element group 324: marked-successors 
    -- CP-element group 324: 	322 
    -- CP-element group 324:  members (3) 
      -- CP-element group 324: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1042_update_completed_
      -- CP-element group 324: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1042_Update/ack
      -- CP-element group 324: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1042_Update/$exit
      -- 
    ack_2207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 324_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend214_exec_guard_965_delayed_1_0_1040_inst_ack_1, ack => zeropad3D_CP_676_elements(324)); -- 
    -- CP-element group 325:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	256 
    -- CP-element group 325: 	264 
    -- CP-element group 325: 	268 
    -- CP-element group 325: 	272 
    -- CP-element group 325: marked-predecessors 
    -- CP-element group 325: 	327 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	327 
    -- CP-element group 325:  members (3) 
      -- CP-element group 325: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1051_Sample/req
      -- CP-element group 325: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1051_Sample/$entry
      -- CP-element group 325: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1051_sample_start_
      -- 
    req_2215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(325), ack => W_ifx_xend214_exec_guard_971_delayed_1_0_1049_inst_req_0); -- 
    zeropad3D_cp_element_group_325: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_325"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(256) & zeropad3D_CP_676_elements(264) & zeropad3D_CP_676_elements(268) & zeropad3D_CP_676_elements(272) & zeropad3D_CP_676_elements(327);
      gj_zeropad3D_cp_element_group_325 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(325), clk => clk, reset => reset); --
    end block;
    -- CP-element group 326:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: marked-predecessors 
    -- CP-element group 326: 	328 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	328 
    -- CP-element group 326:  members (3) 
      -- CP-element group 326: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1051_Update/req
      -- CP-element group 326: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1051_Update/$entry
      -- CP-element group 326: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1051_update_start_
      -- 
    req_2220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(326), ack => W_ifx_xend214_exec_guard_971_delayed_1_0_1049_inst_req_1); -- 
    zeropad3D_cp_element_group_326: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_326"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad3D_CP_676_elements(328);
      gj_zeropad3D_cp_element_group_326 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(326), clk => clk, reset => reset); --
    end block;
    -- CP-element group 327:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	325 
    -- CP-element group 327: successors 
    -- CP-element group 327: marked-successors 
    -- CP-element group 327: 	325 
    -- CP-element group 327: 	254 
    -- CP-element group 327: 	262 
    -- CP-element group 327: 	266 
    -- CP-element group 327: 	270 
    -- CP-element group 327:  members (3) 
      -- CP-element group 327: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1051_Sample/ack
      -- CP-element group 327: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1051_Sample/$exit
      -- CP-element group 327: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1051_sample_completed_
      -- 
    ack_2216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 327_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend214_exec_guard_971_delayed_1_0_1049_inst_ack_0, ack => zeropad3D_CP_676_elements(327)); -- 
    -- CP-element group 328:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	326 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	496 
    -- CP-element group 328: marked-successors 
    -- CP-element group 328: 	326 
    -- CP-element group 328:  members (3) 
      -- CP-element group 328: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1051_Update/ack
      -- CP-element group 328: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1051_Update/$exit
      -- CP-element group 328: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1051_update_completed_
      -- 
    ack_2221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 328_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend214_exec_guard_971_delayed_1_0_1049_inst_ack_1, ack => zeropad3D_CP_676_elements(328)); -- 
    -- CP-element group 329:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	256 
    -- CP-element group 329: 	264 
    -- CP-element group 329: 	268 
    -- CP-element group 329: 	272 
    -- CP-element group 329: marked-predecessors 
    -- CP-element group 329: 	331 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	331 
    -- CP-element group 329:  members (3) 
      -- CP-element group 329: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1061_Sample/$entry
      -- CP-element group 329: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1061_Sample/req
      -- CP-element group 329: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1061_sample_start_
      -- 
    req_2229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(329), ack => W_ifx_xend214_exec_guard_978_delayed_1_0_1059_inst_req_0); -- 
    zeropad3D_cp_element_group_329: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_329"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(256) & zeropad3D_CP_676_elements(264) & zeropad3D_CP_676_elements(268) & zeropad3D_CP_676_elements(272) & zeropad3D_CP_676_elements(331);
      gj_zeropad3D_cp_element_group_329 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(329), clk => clk, reset => reset); --
    end block;
    -- CP-element group 330:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: marked-predecessors 
    -- CP-element group 330: 	332 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	332 
    -- CP-element group 330:  members (3) 
      -- CP-element group 330: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1061_Update/$entry
      -- CP-element group 330: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1061_update_start_
      -- CP-element group 330: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1061_Update/req
      -- 
    req_2234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(330), ack => W_ifx_xend214_exec_guard_978_delayed_1_0_1059_inst_req_1); -- 
    zeropad3D_cp_element_group_330: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_330"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad3D_CP_676_elements(332);
      gj_zeropad3D_cp_element_group_330 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(330), clk => clk, reset => reset); --
    end block;
    -- CP-element group 331:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	329 
    -- CP-element group 331: successors 
    -- CP-element group 331: marked-successors 
    -- CP-element group 331: 	329 
    -- CP-element group 331: 	254 
    -- CP-element group 331: 	262 
    -- CP-element group 331: 	266 
    -- CP-element group 331: 	270 
    -- CP-element group 331:  members (3) 
      -- CP-element group 331: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1061_Sample/ack
      -- CP-element group 331: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1061_Sample/$exit
      -- CP-element group 331: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1061_sample_completed_
      -- 
    ack_2230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 331_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend214_exec_guard_978_delayed_1_0_1059_inst_ack_0, ack => zeropad3D_CP_676_elements(331)); -- 
    -- CP-element group 332:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	330 
    -- CP-element group 332: successors 
    -- CP-element group 332: 	496 
    -- CP-element group 332: marked-successors 
    -- CP-element group 332: 	330 
    -- CP-element group 332:  members (3) 
      -- CP-element group 332: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1061_Update/$exit
      -- CP-element group 332: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1061_update_completed_
      -- CP-element group 332: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1061_Update/ack
      -- 
    ack_2235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend214_exec_guard_978_delayed_1_0_1059_inst_ack_1, ack => zeropad3D_CP_676_elements(332)); -- 
    -- CP-element group 333:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	134 
    -- CP-element group 333: marked-predecessors 
    -- CP-element group 333: 	335 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	335 
    -- CP-element group 333:  members (3) 
      -- CP-element group 333: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1064_Sample/$entry
      -- CP-element group 333: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1064_Sample/rr
      -- CP-element group 333: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1064_sample_start_
      -- 
    rr_2243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(333), ack => type_cast_1064_inst_req_0); -- 
    zeropad3D_cp_element_group_333: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_333"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(134) & zeropad3D_CP_676_elements(335);
      gj_zeropad3D_cp_element_group_333 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(333), clk => clk, reset => reset); --
    end block;
    -- CP-element group 334:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: marked-predecessors 
    -- CP-element group 334: 	336 
    -- CP-element group 334: 	355 
    -- CP-element group 334: 	359 
    -- CP-element group 334: 	363 
    -- CP-element group 334: 	367 
    -- CP-element group 334: 	375 
    -- CP-element group 334: 	379 
    -- CP-element group 334: 	383 
    -- CP-element group 334: 	387 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	336 
    -- CP-element group 334:  members (3) 
      -- CP-element group 334: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1064_Update/$entry
      -- CP-element group 334: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1064_update_start_
      -- CP-element group 334: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1064_Update/cr
      -- 
    cr_2248_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2248_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(334), ack => type_cast_1064_inst_req_1); -- 
    zeropad3D_cp_element_group_334: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_334"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(336) & zeropad3D_CP_676_elements(355) & zeropad3D_CP_676_elements(359) & zeropad3D_CP_676_elements(363) & zeropad3D_CP_676_elements(367) & zeropad3D_CP_676_elements(375) & zeropad3D_CP_676_elements(379) & zeropad3D_CP_676_elements(383) & zeropad3D_CP_676_elements(387);
      gj_zeropad3D_cp_element_group_334 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(334), clk => clk, reset => reset); --
    end block;
    -- CP-element group 335:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	333 
    -- CP-element group 335: successors 
    -- CP-element group 335: marked-successors 
    -- CP-element group 335: 	333 
    -- CP-element group 335:  members (3) 
      -- CP-element group 335: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1064_Sample/$exit
      -- CP-element group 335: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1064_Sample/ra
      -- CP-element group 335: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1064_sample_completed_
      -- 
    ra_2244_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 335_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1064_inst_ack_0, ack => zeropad3D_CP_676_elements(335)); -- 
    -- CP-element group 336:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	334 
    -- CP-element group 336: successors 
    -- CP-element group 336: 	353 
    -- CP-element group 336: 	357 
    -- CP-element group 336: 	361 
    -- CP-element group 336: 	365 
    -- CP-element group 336: 	373 
    -- CP-element group 336: 	377 
    -- CP-element group 336: 	381 
    -- CP-element group 336: 	385 
    -- CP-element group 336: marked-successors 
    -- CP-element group 336: 	334 
    -- CP-element group 336:  members (3) 
      -- CP-element group 336: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1064_Update/$exit
      -- CP-element group 336: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1064_update_completed_
      -- CP-element group 336: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1064_Update/ca
      -- 
    ca_2249_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1064_inst_ack_1, ack => zeropad3D_CP_676_elements(336)); -- 
    -- CP-element group 337:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	256 
    -- CP-element group 337: 	264 
    -- CP-element group 337: 	268 
    -- CP-element group 337: 	272 
    -- CP-element group 337: marked-predecessors 
    -- CP-element group 337: 	339 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	339 
    -- CP-element group 337:  members (3) 
      -- CP-element group 337: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1075_Sample/$entry
      -- CP-element group 337: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1075_sample_start_
      -- CP-element group 337: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1075_Sample/req
      -- 
    req_2257_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2257_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(337), ack => W_ifx_xend214_exec_guard_986_delayed_1_0_1073_inst_req_0); -- 
    zeropad3D_cp_element_group_337: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_337"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(256) & zeropad3D_CP_676_elements(264) & zeropad3D_CP_676_elements(268) & zeropad3D_CP_676_elements(272) & zeropad3D_CP_676_elements(339);
      gj_zeropad3D_cp_element_group_337 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(337), clk => clk, reset => reset); --
    end block;
    -- CP-element group 338:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: marked-predecessors 
    -- CP-element group 338: 	340 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	340 
    -- CP-element group 338:  members (3) 
      -- CP-element group 338: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1075_update_start_
      -- CP-element group 338: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1075_Update/req
      -- CP-element group 338: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1075_Update/$entry
      -- 
    req_2262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(338), ack => W_ifx_xend214_exec_guard_986_delayed_1_0_1073_inst_req_1); -- 
    zeropad3D_cp_element_group_338: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_338"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad3D_CP_676_elements(340);
      gj_zeropad3D_cp_element_group_338 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(338), clk => clk, reset => reset); --
    end block;
    -- CP-element group 339:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	337 
    -- CP-element group 339: successors 
    -- CP-element group 339: marked-successors 
    -- CP-element group 339: 	337 
    -- CP-element group 339: 	254 
    -- CP-element group 339: 	262 
    -- CP-element group 339: 	266 
    -- CP-element group 339: 	270 
    -- CP-element group 339:  members (3) 
      -- CP-element group 339: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1075_Sample/$exit
      -- CP-element group 339: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1075_sample_completed_
      -- CP-element group 339: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1075_Sample/ack
      -- 
    ack_2258_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 339_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend214_exec_guard_986_delayed_1_0_1073_inst_ack_0, ack => zeropad3D_CP_676_elements(339)); -- 
    -- CP-element group 340:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	338 
    -- CP-element group 340: successors 
    -- CP-element group 340: 	496 
    -- CP-element group 340: marked-successors 
    -- CP-element group 340: 	338 
    -- CP-element group 340:  members (3) 
      -- CP-element group 340: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1075_update_completed_
      -- CP-element group 340: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1075_Update/ack
      -- CP-element group 340: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1075_Update/$exit
      -- 
    ack_2263_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend214_exec_guard_986_delayed_1_0_1073_inst_ack_1, ack => zeropad3D_CP_676_elements(340)); -- 
    -- CP-element group 341:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	256 
    -- CP-element group 341: 	264 
    -- CP-element group 341: 	268 
    -- CP-element group 341: 	272 
    -- CP-element group 341: marked-predecessors 
    -- CP-element group 341: 	343 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	343 
    -- CP-element group 341:  members (3) 
      -- CP-element group 341: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1084_sample_start_
      -- CP-element group 341: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1084_Sample/req
      -- CP-element group 341: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1084_Sample/$entry
      -- 
    req_2271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(341), ack => W_ifx_xend214_exec_guard_993_delayed_1_0_1082_inst_req_0); -- 
    zeropad3D_cp_element_group_341: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_341"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(256) & zeropad3D_CP_676_elements(264) & zeropad3D_CP_676_elements(268) & zeropad3D_CP_676_elements(272) & zeropad3D_CP_676_elements(343);
      gj_zeropad3D_cp_element_group_341 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(341), clk => clk, reset => reset); --
    end block;
    -- CP-element group 342:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: marked-predecessors 
    -- CP-element group 342: 	344 
    -- CP-element group 342: 	355 
    -- CP-element group 342: 	359 
    -- CP-element group 342: 	363 
    -- CP-element group 342: 	367 
    -- CP-element group 342: 	375 
    -- CP-element group 342: 	379 
    -- CP-element group 342: 	383 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	344 
    -- CP-element group 342:  members (3) 
      -- CP-element group 342: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1084_Update/$entry
      -- CP-element group 342: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1084_Update/req
      -- CP-element group 342: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1084_update_start_
      -- 
    req_2276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(342), ack => W_ifx_xend214_exec_guard_993_delayed_1_0_1082_inst_req_1); -- 
    zeropad3D_cp_element_group_342: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_342"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(344) & zeropad3D_CP_676_elements(355) & zeropad3D_CP_676_elements(359) & zeropad3D_CP_676_elements(363) & zeropad3D_CP_676_elements(367) & zeropad3D_CP_676_elements(375) & zeropad3D_CP_676_elements(379) & zeropad3D_CP_676_elements(383);
      gj_zeropad3D_cp_element_group_342 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(342), clk => clk, reset => reset); --
    end block;
    -- CP-element group 343:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	341 
    -- CP-element group 343: successors 
    -- CP-element group 343: marked-successors 
    -- CP-element group 343: 	341 
    -- CP-element group 343: 	254 
    -- CP-element group 343: 	262 
    -- CP-element group 343: 	266 
    -- CP-element group 343: 	270 
    -- CP-element group 343:  members (3) 
      -- CP-element group 343: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1084_Sample/$exit
      -- CP-element group 343: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1084_sample_completed_
      -- CP-element group 343: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1084_Sample/ack
      -- 
    ack_2272_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 343_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend214_exec_guard_993_delayed_1_0_1082_inst_ack_0, ack => zeropad3D_CP_676_elements(343)); -- 
    -- CP-element group 344:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	342 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	353 
    -- CP-element group 344: 	357 
    -- CP-element group 344: 	361 
    -- CP-element group 344: 	365 
    -- CP-element group 344: 	373 
    -- CP-element group 344: 	377 
    -- CP-element group 344: 	381 
    -- CP-element group 344: marked-successors 
    -- CP-element group 344: 	342 
    -- CP-element group 344:  members (3) 
      -- CP-element group 344: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1084_update_completed_
      -- CP-element group 344: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1084_Update/$exit
      -- CP-element group 344: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1084_Update/ack
      -- 
    ack_2277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 344_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend214_exec_guard_993_delayed_1_0_1082_inst_ack_1, ack => zeropad3D_CP_676_elements(344)); -- 
    -- CP-element group 345:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	256 
    -- CP-element group 345: 	264 
    -- CP-element group 345: 	268 
    -- CP-element group 345: 	272 
    -- CP-element group 345: marked-predecessors 
    -- CP-element group 345: 	347 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	347 
    -- CP-element group 345:  members (3) 
      -- CP-element group 345: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1092_Sample/req
      -- CP-element group 345: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1092_Sample/$entry
      -- CP-element group 345: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1092_sample_start_
      -- 
    req_2285_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2285_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(345), ack => W_ifx_xend214_exec_guard_998_delayed_1_0_1090_inst_req_0); -- 
    zeropad3D_cp_element_group_345: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_345"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(256) & zeropad3D_CP_676_elements(264) & zeropad3D_CP_676_elements(268) & zeropad3D_CP_676_elements(272) & zeropad3D_CP_676_elements(347);
      gj_zeropad3D_cp_element_group_345 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(345), clk => clk, reset => reset); --
    end block;
    -- CP-element group 346:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: marked-predecessors 
    -- CP-element group 346: 	348 
    -- CP-element group 346: 	387 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	348 
    -- CP-element group 346:  members (3) 
      -- CP-element group 346: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1092_Update/req
      -- CP-element group 346: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1092_Update/$entry
      -- CP-element group 346: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1092_update_start_
      -- 
    req_2290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(346), ack => W_ifx_xend214_exec_guard_998_delayed_1_0_1090_inst_req_1); -- 
    zeropad3D_cp_element_group_346: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_346"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(348) & zeropad3D_CP_676_elements(387);
      gj_zeropad3D_cp_element_group_346 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(346), clk => clk, reset => reset); --
    end block;
    -- CP-element group 347:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	345 
    -- CP-element group 347: successors 
    -- CP-element group 347: marked-successors 
    -- CP-element group 347: 	345 
    -- CP-element group 347: 	254 
    -- CP-element group 347: 	262 
    -- CP-element group 347: 	266 
    -- CP-element group 347: 	270 
    -- CP-element group 347:  members (3) 
      -- CP-element group 347: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1092_Sample/ack
      -- CP-element group 347: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1092_Sample/$exit
      -- CP-element group 347: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1092_sample_completed_
      -- 
    ack_2286_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 347_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend214_exec_guard_998_delayed_1_0_1090_inst_ack_0, ack => zeropad3D_CP_676_elements(347)); -- 
    -- CP-element group 348:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	346 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	385 
    -- CP-element group 348: marked-successors 
    -- CP-element group 348: 	346 
    -- CP-element group 348:  members (3) 
      -- CP-element group 348: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1092_Update/ack
      -- CP-element group 348: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1092_Update/$exit
      -- CP-element group 348: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1092_update_completed_
      -- 
    ack_2291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 348_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend214_exec_guard_998_delayed_1_0_1090_inst_ack_1, ack => zeropad3D_CP_676_elements(348)); -- 
    -- CP-element group 349:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	300 
    -- CP-element group 349: 	304 
    -- CP-element group 349: 	308 
    -- CP-element group 349: 	312 
    -- CP-element group 349: 	256 
    -- CP-element group 349: 	264 
    -- CP-element group 349: 	268 
    -- CP-element group 349: marked-predecessors 
    -- CP-element group 349: 	351 
    -- CP-element group 349: successors 
    -- CP-element group 349: 	351 
    -- CP-element group 349:  members (3) 
      -- CP-element group 349: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1104_Sample/req
      -- CP-element group 349: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1104_Sample/$entry
      -- CP-element group 349: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1104_sample_start_
      -- 
    req_2299_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2299_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(349), ack => W_jx_x0_1008_delayed_1_0_1102_inst_req_0); -- 
    zeropad3D_cp_element_group_349: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_349"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(300) & zeropad3D_CP_676_elements(304) & zeropad3D_CP_676_elements(308) & zeropad3D_CP_676_elements(312) & zeropad3D_CP_676_elements(256) & zeropad3D_CP_676_elements(264) & zeropad3D_CP_676_elements(268) & zeropad3D_CP_676_elements(351);
      gj_zeropad3D_cp_element_group_349 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(349), clk => clk, reset => reset); --
    end block;
    -- CP-element group 350:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: marked-predecessors 
    -- CP-element group 350: 	352 
    -- CP-element group 350: 	355 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	352 
    -- CP-element group 350:  members (3) 
      -- CP-element group 350: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1104_Update/req
      -- CP-element group 350: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1104_Update/$entry
      -- CP-element group 350: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1104_update_start_
      -- 
    req_2304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(350), ack => W_jx_x0_1008_delayed_1_0_1102_inst_req_1); -- 
    zeropad3D_cp_element_group_350: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_350"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(352) & zeropad3D_CP_676_elements(355);
      gj_zeropad3D_cp_element_group_350 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(350), clk => clk, reset => reset); --
    end block;
    -- CP-element group 351:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	349 
    -- CP-element group 351: successors 
    -- CP-element group 351: marked-successors 
    -- CP-element group 351: 	349 
    -- CP-element group 351: 	298 
    -- CP-element group 351: 	302 
    -- CP-element group 351: 	306 
    -- CP-element group 351: 	310 
    -- CP-element group 351: 	254 
    -- CP-element group 351: 	262 
    -- CP-element group 351: 	266 
    -- CP-element group 351:  members (3) 
      -- CP-element group 351: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1104_Sample/ack
      -- CP-element group 351: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1104_Sample/$exit
      -- CP-element group 351: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1104_sample_completed_
      -- 
    ack_2300_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 351_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_jx_x0_1008_delayed_1_0_1102_inst_ack_0, ack => zeropad3D_CP_676_elements(351)); -- 
    -- CP-element group 352:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	350 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	353 
    -- CP-element group 352: marked-successors 
    -- CP-element group 352: 	350 
    -- CP-element group 352:  members (3) 
      -- CP-element group 352: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1104_Update/ack
      -- CP-element group 352: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1104_Update/$exit
      -- CP-element group 352: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1104_update_completed_
      -- 
    ack_2305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_jx_x0_1008_delayed_1_0_1102_inst_ack_1, ack => zeropad3D_CP_676_elements(352)); -- 
    -- CP-element group 353:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	336 
    -- CP-element group 353: 	344 
    -- CP-element group 353: 	352 
    -- CP-element group 353: 	320 
    -- CP-element group 353: marked-predecessors 
    -- CP-element group 353: 	355 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	355 
    -- CP-element group 353:  members (3) 
      -- CP-element group 353: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1108_Sample/$entry
      -- CP-element group 353: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1108_sample_start_
      -- CP-element group 353: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1108_Sample/rr
      -- 
    rr_2313_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2313_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(353), ack => type_cast_1108_inst_req_0); -- 
    zeropad3D_cp_element_group_353: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_353"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(336) & zeropad3D_CP_676_elements(344) & zeropad3D_CP_676_elements(352) & zeropad3D_CP_676_elements(320) & zeropad3D_CP_676_elements(355);
      gj_zeropad3D_cp_element_group_353 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(353), clk => clk, reset => reset); --
    end block;
    -- CP-element group 354:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: marked-predecessors 
    -- CP-element group 354: 	356 
    -- CP-element group 354: 	395 
    -- CP-element group 354: 	399 
    -- CP-element group 354: 	403 
    -- CP-element group 354: 	426 
    -- CP-element group 354: 	430 
    -- CP-element group 354: 	434 
    -- CP-element group 354: 	449 
    -- CP-element group 354: 	461 
    -- CP-element group 354: 	465 
    -- CP-element group 354: 	469 
    -- CP-element group 354: 	484 
    -- CP-element group 354: successors 
    -- CP-element group 354: 	356 
    -- CP-element group 354:  members (3) 
      -- CP-element group 354: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1108_Update/$entry
      -- CP-element group 354: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1108_Update/cr
      -- CP-element group 354: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1108_update_start_
      -- 
    cr_2318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(354), ack => type_cast_1108_inst_req_1); -- 
    zeropad3D_cp_element_group_354: block -- 
      constant place_capacities: IntegerArray(0 to 11) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_markings: IntegerArray(0 to 11)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_delays: IntegerArray(0 to 11) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_354"; 
      signal preds: BooleanArray(1 to 12); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(356) & zeropad3D_CP_676_elements(395) & zeropad3D_CP_676_elements(399) & zeropad3D_CP_676_elements(403) & zeropad3D_CP_676_elements(426) & zeropad3D_CP_676_elements(430) & zeropad3D_CP_676_elements(434) & zeropad3D_CP_676_elements(449) & zeropad3D_CP_676_elements(461) & zeropad3D_CP_676_elements(465) & zeropad3D_CP_676_elements(469) & zeropad3D_CP_676_elements(484);
      gj_zeropad3D_cp_element_group_354 : generic_join generic map(name => joinName, number_of_predecessors => 12, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(354), clk => clk, reset => reset); --
    end block;
    -- CP-element group 355:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	353 
    -- CP-element group 355: successors 
    -- CP-element group 355: marked-successors 
    -- CP-element group 355: 	334 
    -- CP-element group 355: 	342 
    -- CP-element group 355: 	350 
    -- CP-element group 355: 	353 
    -- CP-element group 355: 	318 
    -- CP-element group 355:  members (3) 
      -- CP-element group 355: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1108_Sample/ra
      -- CP-element group 355: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1108_sample_completed_
      -- CP-element group 355: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1108_Sample/$exit
      -- 
    ra_2314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 355_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1108_inst_ack_0, ack => zeropad3D_CP_676_elements(355)); -- 
    -- CP-element group 356:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	354 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	393 
    -- CP-element group 356: 	397 
    -- CP-element group 356: 	401 
    -- CP-element group 356: 	424 
    -- CP-element group 356: 	428 
    -- CP-element group 356: 	432 
    -- CP-element group 356: 	447 
    -- CP-element group 356: 	459 
    -- CP-element group 356: 	463 
    -- CP-element group 356: 	467 
    -- CP-element group 356: 	482 
    -- CP-element group 356: marked-successors 
    -- CP-element group 356: 	354 
    -- CP-element group 356:  members (3) 
      -- CP-element group 356: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1108_update_completed_
      -- CP-element group 356: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1108_Update/ca
      -- CP-element group 356: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1108_Update/$exit
      -- 
    ca_2319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 356_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1108_inst_ack_1, ack => zeropad3D_CP_676_elements(356)); -- 
    -- CP-element group 357:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	336 
    -- CP-element group 357: 	344 
    -- CP-element group 357: 	320 
    -- CP-element group 357: marked-predecessors 
    -- CP-element group 357: 	359 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	359 
    -- CP-element group 357:  members (3) 
      -- CP-element group 357: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1112_sample_start_
      -- CP-element group 357: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1112_Sample/req
      -- CP-element group 357: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1112_Sample/$entry
      -- 
    req_2327_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2327_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(357), ack => W_lorx_xlhsx_xfalse269_exec_guard_1011_delayed_1_0_1110_inst_req_0); -- 
    zeropad3D_cp_element_group_357: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_357"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(336) & zeropad3D_CP_676_elements(344) & zeropad3D_CP_676_elements(320) & zeropad3D_CP_676_elements(359);
      gj_zeropad3D_cp_element_group_357 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(357), clk => clk, reset => reset); --
    end block;
    -- CP-element group 358:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: marked-predecessors 
    -- CP-element group 358: 	360 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	360 
    -- CP-element group 358:  members (3) 
      -- CP-element group 358: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1112_update_start_
      -- CP-element group 358: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1112_Update/req
      -- CP-element group 358: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1112_Update/$entry
      -- 
    req_2332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(358), ack => W_lorx_xlhsx_xfalse269_exec_guard_1011_delayed_1_0_1110_inst_req_1); -- 
    zeropad3D_cp_element_group_358: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_358"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad3D_CP_676_elements(360);
      gj_zeropad3D_cp_element_group_358 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(358), clk => clk, reset => reset); --
    end block;
    -- CP-element group 359:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	357 
    -- CP-element group 359: successors 
    -- CP-element group 359: marked-successors 
    -- CP-element group 359: 	334 
    -- CP-element group 359: 	342 
    -- CP-element group 359: 	357 
    -- CP-element group 359: 	318 
    -- CP-element group 359:  members (3) 
      -- CP-element group 359: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1112_sample_completed_
      -- CP-element group 359: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1112_Sample/ack
      -- CP-element group 359: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1112_Sample/$exit
      -- 
    ack_2328_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 359_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_lorx_xlhsx_xfalse269_exec_guard_1011_delayed_1_0_1110_inst_ack_0, ack => zeropad3D_CP_676_elements(359)); -- 
    -- CP-element group 360:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	358 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	496 
    -- CP-element group 360: marked-successors 
    -- CP-element group 360: 	358 
    -- CP-element group 360:  members (3) 
      -- CP-element group 360: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1112_update_completed_
      -- CP-element group 360: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1112_Update/ack
      -- CP-element group 360: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1112_Update/$exit
      -- 
    ack_2333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 360_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_lorx_xlhsx_xfalse269_exec_guard_1011_delayed_1_0_1110_inst_ack_1, ack => zeropad3D_CP_676_elements(360)); -- 
    -- CP-element group 361:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	336 
    -- CP-element group 361: 	344 
    -- CP-element group 361: 	320 
    -- CP-element group 361: marked-predecessors 
    -- CP-element group 361: 	363 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	363 
    -- CP-element group 361:  members (3) 
      -- CP-element group 361: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1121_Sample/req
      -- CP-element group 361: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1121_Sample/$entry
      -- CP-element group 361: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1121_sample_start_
      -- 
    req_2341_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2341_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(361), ack => W_lorx_xlhsx_xfalse269_exec_guard_1017_delayed_1_0_1119_inst_req_0); -- 
    zeropad3D_cp_element_group_361: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_361"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(336) & zeropad3D_CP_676_elements(344) & zeropad3D_CP_676_elements(320) & zeropad3D_CP_676_elements(363);
      gj_zeropad3D_cp_element_group_361 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(361), clk => clk, reset => reset); --
    end block;
    -- CP-element group 362:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: marked-predecessors 
    -- CP-element group 362: 	364 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	364 
    -- CP-element group 362:  members (3) 
      -- CP-element group 362: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1121_Update/req
      -- CP-element group 362: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1121_Update/$entry
      -- CP-element group 362: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1121_update_start_
      -- 
    req_2346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(362), ack => W_lorx_xlhsx_xfalse269_exec_guard_1017_delayed_1_0_1119_inst_req_1); -- 
    zeropad3D_cp_element_group_362: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_362"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad3D_CP_676_elements(364);
      gj_zeropad3D_cp_element_group_362 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(362), clk => clk, reset => reset); --
    end block;
    -- CP-element group 363:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	361 
    -- CP-element group 363: successors 
    -- CP-element group 363: marked-successors 
    -- CP-element group 363: 	334 
    -- CP-element group 363: 	342 
    -- CP-element group 363: 	361 
    -- CP-element group 363: 	318 
    -- CP-element group 363:  members (3) 
      -- CP-element group 363: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1121_Sample/ack
      -- CP-element group 363: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1121_Sample/$exit
      -- CP-element group 363: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1121_sample_completed_
      -- 
    ack_2342_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 363_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_lorx_xlhsx_xfalse269_exec_guard_1017_delayed_1_0_1119_inst_ack_0, ack => zeropad3D_CP_676_elements(363)); -- 
    -- CP-element group 364:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	362 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	496 
    -- CP-element group 364: marked-successors 
    -- CP-element group 364: 	362 
    -- CP-element group 364:  members (3) 
      -- CP-element group 364: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1121_Update/ack
      -- CP-element group 364: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1121_Update/$exit
      -- CP-element group 364: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1121_update_completed_
      -- 
    ack_2347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 364_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_lorx_xlhsx_xfalse269_exec_guard_1017_delayed_1_0_1119_inst_ack_1, ack => zeropad3D_CP_676_elements(364)); -- 
    -- CP-element group 365:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	336 
    -- CP-element group 365: 	344 
    -- CP-element group 365: 	320 
    -- CP-element group 365: marked-predecessors 
    -- CP-element group 365: 	367 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	367 
    -- CP-element group 365:  members (3) 
      -- CP-element group 365: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1131_sample_start_
      -- CP-element group 365: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1131_Sample/req
      -- CP-element group 365: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1131_Sample/$entry
      -- 
    req_2355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(365), ack => W_lorx_xlhsx_xfalse269_exec_guard_1024_delayed_1_0_1129_inst_req_0); -- 
    zeropad3D_cp_element_group_365: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_365"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(336) & zeropad3D_CP_676_elements(344) & zeropad3D_CP_676_elements(320) & zeropad3D_CP_676_elements(367);
      gj_zeropad3D_cp_element_group_365 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(365), clk => clk, reset => reset); --
    end block;
    -- CP-element group 366:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: marked-predecessors 
    -- CP-element group 366: 	368 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	368 
    -- CP-element group 366:  members (3) 
      -- CP-element group 366: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1131_Update/req
      -- CP-element group 366: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1131_Update/$entry
      -- CP-element group 366: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1131_update_start_
      -- 
    req_2360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(366), ack => W_lorx_xlhsx_xfalse269_exec_guard_1024_delayed_1_0_1129_inst_req_1); -- 
    zeropad3D_cp_element_group_366: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_366"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad3D_CP_676_elements(368);
      gj_zeropad3D_cp_element_group_366 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(366), clk => clk, reset => reset); --
    end block;
    -- CP-element group 367:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	365 
    -- CP-element group 367: successors 
    -- CP-element group 367: marked-successors 
    -- CP-element group 367: 	334 
    -- CP-element group 367: 	342 
    -- CP-element group 367: 	365 
    -- CP-element group 367: 	318 
    -- CP-element group 367:  members (3) 
      -- CP-element group 367: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1131_Sample/ack
      -- CP-element group 367: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1131_Sample/$exit
      -- CP-element group 367: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1131_sample_completed_
      -- 
    ack_2356_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 367_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_lorx_xlhsx_xfalse269_exec_guard_1024_delayed_1_0_1129_inst_ack_0, ack => zeropad3D_CP_676_elements(367)); -- 
    -- CP-element group 368:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	366 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	496 
    -- CP-element group 368: marked-successors 
    -- CP-element group 368: 	366 
    -- CP-element group 368:  members (3) 
      -- CP-element group 368: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1131_Update/ack
      -- CP-element group 368: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1131_Update/$exit
      -- CP-element group 368: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1131_update_completed_
      -- 
    ack_2361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 368_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_lorx_xlhsx_xfalse269_exec_guard_1024_delayed_1_0_1129_inst_ack_1, ack => zeropad3D_CP_676_elements(368)); -- 
    -- CP-element group 369:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	134 
    -- CP-element group 369: marked-predecessors 
    -- CP-element group 369: 	371 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	371 
    -- CP-element group 369:  members (3) 
      -- CP-element group 369: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1134_sample_start_
      -- CP-element group 369: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1134_Sample/rr
      -- CP-element group 369: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1134_Sample/$entry
      -- 
    rr_2369_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2369_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(369), ack => type_cast_1134_inst_req_0); -- 
    zeropad3D_cp_element_group_369: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_369"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(134) & zeropad3D_CP_676_elements(371);
      gj_zeropad3D_cp_element_group_369 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(369), clk => clk, reset => reset); --
    end block;
    -- CP-element group 370:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: marked-predecessors 
    -- CP-element group 370: 	372 
    -- CP-element group 370: 	395 
    -- CP-element group 370: 	399 
    -- CP-element group 370: 	403 
    -- CP-element group 370: 	426 
    -- CP-element group 370: 	430 
    -- CP-element group 370: 	434 
    -- CP-element group 370: 	449 
    -- CP-element group 370: 	461 
    -- CP-element group 370: 	465 
    -- CP-element group 370: 	469 
    -- CP-element group 370: 	484 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	372 
    -- CP-element group 370:  members (3) 
      -- CP-element group 370: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1134_update_start_
      -- CP-element group 370: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1134_Update/$entry
      -- CP-element group 370: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1134_Update/cr
      -- 
    cr_2374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(370), ack => type_cast_1134_inst_req_1); -- 
    zeropad3D_cp_element_group_370: block -- 
      constant place_capacities: IntegerArray(0 to 11) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_markings: IntegerArray(0 to 11)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_delays: IntegerArray(0 to 11) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_370"; 
      signal preds: BooleanArray(1 to 12); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(372) & zeropad3D_CP_676_elements(395) & zeropad3D_CP_676_elements(399) & zeropad3D_CP_676_elements(403) & zeropad3D_CP_676_elements(426) & zeropad3D_CP_676_elements(430) & zeropad3D_CP_676_elements(434) & zeropad3D_CP_676_elements(449) & zeropad3D_CP_676_elements(461) & zeropad3D_CP_676_elements(465) & zeropad3D_CP_676_elements(469) & zeropad3D_CP_676_elements(484);
      gj_zeropad3D_cp_element_group_370 : generic_join generic map(name => joinName, number_of_predecessors => 12, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(370), clk => clk, reset => reset); --
    end block;
    -- CP-element group 371:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	369 
    -- CP-element group 371: successors 
    -- CP-element group 371: marked-successors 
    -- CP-element group 371: 	369 
    -- CP-element group 371:  members (3) 
      -- CP-element group 371: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1134_sample_completed_
      -- CP-element group 371: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1134_Sample/ra
      -- CP-element group 371: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1134_Sample/$exit
      -- 
    ra_2370_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 371_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1134_inst_ack_0, ack => zeropad3D_CP_676_elements(371)); -- 
    -- CP-element group 372:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	370 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	393 
    -- CP-element group 372: 	397 
    -- CP-element group 372: 	401 
    -- CP-element group 372: 	424 
    -- CP-element group 372: 	428 
    -- CP-element group 372: 	432 
    -- CP-element group 372: 	447 
    -- CP-element group 372: 	459 
    -- CP-element group 372: 	463 
    -- CP-element group 372: 	467 
    -- CP-element group 372: 	482 
    -- CP-element group 372: marked-successors 
    -- CP-element group 372: 	370 
    -- CP-element group 372:  members (3) 
      -- CP-element group 372: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1134_update_completed_
      -- CP-element group 372: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1134_Update/$exit
      -- CP-element group 372: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1134_Update/ca
      -- 
    ca_2375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 372_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1134_inst_ack_1, ack => zeropad3D_CP_676_elements(372)); -- 
    -- CP-element group 373:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	336 
    -- CP-element group 373: 	344 
    -- CP-element group 373: 	320 
    -- CP-element group 373: marked-predecessors 
    -- CP-element group 373: 	375 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	375 
    -- CP-element group 373:  members (3) 
      -- CP-element group 373: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1145_sample_start_
      -- CP-element group 373: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1145_Sample/req
      -- CP-element group 373: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1145_Sample/$entry
      -- 
    req_2383_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2383_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(373), ack => W_lorx_xlhsx_xfalse269_exec_guard_1032_delayed_1_0_1143_inst_req_0); -- 
    zeropad3D_cp_element_group_373: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_373"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(336) & zeropad3D_CP_676_elements(344) & zeropad3D_CP_676_elements(320) & zeropad3D_CP_676_elements(375);
      gj_zeropad3D_cp_element_group_373 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(373), clk => clk, reset => reset); --
    end block;
    -- CP-element group 374:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: marked-predecessors 
    -- CP-element group 374: 	376 
    -- CP-element group 374: successors 
    -- CP-element group 374: 	376 
    -- CP-element group 374:  members (3) 
      -- CP-element group 374: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1145_Update/req
      -- CP-element group 374: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1145_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1145_update_start_
      -- 
    req_2388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(374), ack => W_lorx_xlhsx_xfalse269_exec_guard_1032_delayed_1_0_1143_inst_req_1); -- 
    zeropad3D_cp_element_group_374: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_374"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad3D_CP_676_elements(376);
      gj_zeropad3D_cp_element_group_374 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(374), clk => clk, reset => reset); --
    end block;
    -- CP-element group 375:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	373 
    -- CP-element group 375: successors 
    -- CP-element group 375: marked-successors 
    -- CP-element group 375: 	334 
    -- CP-element group 375: 	342 
    -- CP-element group 375: 	318 
    -- CP-element group 375: 	373 
    -- CP-element group 375:  members (3) 
      -- CP-element group 375: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1145_sample_completed_
      -- CP-element group 375: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1145_Sample/ack
      -- CP-element group 375: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1145_Sample/$exit
      -- 
    ack_2384_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 375_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_lorx_xlhsx_xfalse269_exec_guard_1032_delayed_1_0_1143_inst_ack_0, ack => zeropad3D_CP_676_elements(375)); -- 
    -- CP-element group 376:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	374 
    -- CP-element group 376: successors 
    -- CP-element group 376: 	496 
    -- CP-element group 376: marked-successors 
    -- CP-element group 376: 	374 
    -- CP-element group 376:  members (3) 
      -- CP-element group 376: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1145_update_completed_
      -- CP-element group 376: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1145_Update/ack
      -- CP-element group 376: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1145_Update/$exit
      -- 
    ack_2389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 376_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_lorx_xlhsx_xfalse269_exec_guard_1032_delayed_1_0_1143_inst_ack_1, ack => zeropad3D_CP_676_elements(376)); -- 
    -- CP-element group 377:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	336 
    -- CP-element group 377: 	344 
    -- CP-element group 377: 	320 
    -- CP-element group 377: marked-predecessors 
    -- CP-element group 377: 	379 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	379 
    -- CP-element group 377:  members (3) 
      -- CP-element group 377: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1154_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1154_Sample/req
      -- CP-element group 377: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1154_Sample/$entry
      -- 
    req_2397_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2397_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(377), ack => W_lorx_xlhsx_xfalse269_exec_guard_1039_delayed_1_0_1152_inst_req_0); -- 
    zeropad3D_cp_element_group_377: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_377"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(336) & zeropad3D_CP_676_elements(344) & zeropad3D_CP_676_elements(320) & zeropad3D_CP_676_elements(379);
      gj_zeropad3D_cp_element_group_377 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(377), clk => clk, reset => reset); --
    end block;
    -- CP-element group 378:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: marked-predecessors 
    -- CP-element group 378: 	380 
    -- CP-element group 378: 	426 
    -- CP-element group 378: 	430 
    -- CP-element group 378: 	434 
    -- CP-element group 378: 	449 
    -- CP-element group 378: 	461 
    -- CP-element group 378: 	465 
    -- CP-element group 378: 	469 
    -- CP-element group 378: 	484 
    -- CP-element group 378: successors 
    -- CP-element group 378: 	380 
    -- CP-element group 378:  members (3) 
      -- CP-element group 378: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1154_Update/$entry
      -- CP-element group 378: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1154_Update/req
      -- CP-element group 378: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1154_update_start_
      -- 
    req_2402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(378), ack => W_lorx_xlhsx_xfalse269_exec_guard_1039_delayed_1_0_1152_inst_req_1); -- 
    zeropad3D_cp_element_group_378: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_378"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(380) & zeropad3D_CP_676_elements(426) & zeropad3D_CP_676_elements(430) & zeropad3D_CP_676_elements(434) & zeropad3D_CP_676_elements(449) & zeropad3D_CP_676_elements(461) & zeropad3D_CP_676_elements(465) & zeropad3D_CP_676_elements(469) & zeropad3D_CP_676_elements(484);
      gj_zeropad3D_cp_element_group_378 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(378), clk => clk, reset => reset); --
    end block;
    -- CP-element group 379:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	377 
    -- CP-element group 379: successors 
    -- CP-element group 379: marked-successors 
    -- CP-element group 379: 	334 
    -- CP-element group 379: 	342 
    -- CP-element group 379: 	318 
    -- CP-element group 379: 	377 
    -- CP-element group 379:  members (3) 
      -- CP-element group 379: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1154_Sample/ack
      -- CP-element group 379: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1154_Sample/$exit
      -- CP-element group 379: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1154_sample_completed_
      -- 
    ack_2398_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 379_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_lorx_xlhsx_xfalse269_exec_guard_1039_delayed_1_0_1152_inst_ack_0, ack => zeropad3D_CP_676_elements(379)); -- 
    -- CP-element group 380:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	378 
    -- CP-element group 380: successors 
    -- CP-element group 380: 	424 
    -- CP-element group 380: 	428 
    -- CP-element group 380: 	432 
    -- CP-element group 380: 	447 
    -- CP-element group 380: 	459 
    -- CP-element group 380: 	463 
    -- CP-element group 380: 	467 
    -- CP-element group 380: 	482 
    -- CP-element group 380: marked-successors 
    -- CP-element group 380: 	378 
    -- CP-element group 380:  members (3) 
      -- CP-element group 380: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1154_Update/ack
      -- CP-element group 380: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1154_Update/$exit
      -- CP-element group 380: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1154_update_completed_
      -- 
    ack_2403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 380_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_lorx_xlhsx_xfalse269_exec_guard_1039_delayed_1_0_1152_inst_ack_1, ack => zeropad3D_CP_676_elements(380)); -- 
    -- CP-element group 381:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	336 
    -- CP-element group 381: 	344 
    -- CP-element group 381: 	320 
    -- CP-element group 381: marked-predecessors 
    -- CP-element group 381: 	383 
    -- CP-element group 381: successors 
    -- CP-element group 381: 	383 
    -- CP-element group 381:  members (3) 
      -- CP-element group 381: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1162_Sample/req
      -- CP-element group 381: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1162_Sample/$entry
      -- CP-element group 381: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1162_sample_start_
      -- 
    req_2411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(381), ack => W_lorx_xlhsx_xfalse269_exec_guard_1044_delayed_1_0_1160_inst_req_0); -- 
    zeropad3D_cp_element_group_381: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_381"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(336) & zeropad3D_CP_676_elements(344) & zeropad3D_CP_676_elements(320) & zeropad3D_CP_676_elements(383);
      gj_zeropad3D_cp_element_group_381 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(381), clk => clk, reset => reset); --
    end block;
    -- CP-element group 382:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: marked-predecessors 
    -- CP-element group 382: 	384 
    -- CP-element group 382: 	395 
    -- CP-element group 382: 	399 
    -- CP-element group 382: 	403 
    -- CP-element group 382: successors 
    -- CP-element group 382: 	384 
    -- CP-element group 382:  members (3) 
      -- CP-element group 382: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1162_Update/req
      -- CP-element group 382: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1162_Update/$entry
      -- CP-element group 382: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1162_update_start_
      -- 
    req_2416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(382), ack => W_lorx_xlhsx_xfalse269_exec_guard_1044_delayed_1_0_1160_inst_req_1); -- 
    zeropad3D_cp_element_group_382: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_382"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(384) & zeropad3D_CP_676_elements(395) & zeropad3D_CP_676_elements(399) & zeropad3D_CP_676_elements(403);
      gj_zeropad3D_cp_element_group_382 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(382), clk => clk, reset => reset); --
    end block;
    -- CP-element group 383:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	381 
    -- CP-element group 383: successors 
    -- CP-element group 383: marked-successors 
    -- CP-element group 383: 	334 
    -- CP-element group 383: 	342 
    -- CP-element group 383: 	318 
    -- CP-element group 383: 	381 
    -- CP-element group 383:  members (3) 
      -- CP-element group 383: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1162_Sample/ack
      -- CP-element group 383: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1162_Sample/$exit
      -- CP-element group 383: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1162_sample_completed_
      -- 
    ack_2412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 383_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_lorx_xlhsx_xfalse269_exec_guard_1044_delayed_1_0_1160_inst_ack_0, ack => zeropad3D_CP_676_elements(383)); -- 
    -- CP-element group 384:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	382 
    -- CP-element group 384: successors 
    -- CP-element group 384: 	393 
    -- CP-element group 384: 	397 
    -- CP-element group 384: 	401 
    -- CP-element group 384: marked-successors 
    -- CP-element group 384: 	382 
    -- CP-element group 384:  members (3) 
      -- CP-element group 384: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1162_Update/ack
      -- CP-element group 384: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1162_Update/$exit
      -- CP-element group 384: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1162_update_completed_
      -- 
    ack_2417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 384_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_lorx_xlhsx_xfalse269_exec_guard_1044_delayed_1_0_1160_inst_ack_1, ack => zeropad3D_CP_676_elements(384)); -- 
    -- CP-element group 385:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	336 
    -- CP-element group 385: 	348 
    -- CP-element group 385: 	320 
    -- CP-element group 385: marked-predecessors 
    -- CP-element group 385: 	387 
    -- CP-element group 385: successors 
    -- CP-element group 385: 	387 
    -- CP-element group 385:  members (3) 
      -- CP-element group 385: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1171_sample_start_
      -- CP-element group 385: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1171_Sample/req
      -- CP-element group 385: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1171_Sample/$entry
      -- 
    req_2425_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2425_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(385), ack => W_ifx_xend214_ifx_xthen286_taken_1050_delayed_1_0_1169_inst_req_0); -- 
    zeropad3D_cp_element_group_385: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_385"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(336) & zeropad3D_CP_676_elements(348) & zeropad3D_CP_676_elements(320) & zeropad3D_CP_676_elements(387);
      gj_zeropad3D_cp_element_group_385 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(385), clk => clk, reset => reset); --
    end block;
    -- CP-element group 386:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: marked-predecessors 
    -- CP-element group 386: 	388 
    -- CP-element group 386: 	395 
    -- CP-element group 386: 	399 
    -- CP-element group 386: 	403 
    -- CP-element group 386: successors 
    -- CP-element group 386: 	388 
    -- CP-element group 386:  members (3) 
      -- CP-element group 386: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1171_update_start_
      -- CP-element group 386: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1171_Update/req
      -- CP-element group 386: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1171_Update/$entry
      -- 
    req_2430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(386), ack => W_ifx_xend214_ifx_xthen286_taken_1050_delayed_1_0_1169_inst_req_1); -- 
    zeropad3D_cp_element_group_386: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_386"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(388) & zeropad3D_CP_676_elements(395) & zeropad3D_CP_676_elements(399) & zeropad3D_CP_676_elements(403);
      gj_zeropad3D_cp_element_group_386 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(386), clk => clk, reset => reset); --
    end block;
    -- CP-element group 387:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	385 
    -- CP-element group 387: successors 
    -- CP-element group 387: marked-successors 
    -- CP-element group 387: 	334 
    -- CP-element group 387: 	346 
    -- CP-element group 387: 	318 
    -- CP-element group 387: 	385 
    -- CP-element group 387:  members (3) 
      -- CP-element group 387: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1171_Sample/ack
      -- CP-element group 387: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1171_Sample/$exit
      -- CP-element group 387: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1171_sample_completed_
      -- 
    ack_2426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 387_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend214_ifx_xthen286_taken_1050_delayed_1_0_1169_inst_ack_0, ack => zeropad3D_CP_676_elements(387)); -- 
    -- CP-element group 388:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: 	386 
    -- CP-element group 388: successors 
    -- CP-element group 388: 	393 
    -- CP-element group 388: 	397 
    -- CP-element group 388: 	401 
    -- CP-element group 388: marked-successors 
    -- CP-element group 388: 	386 
    -- CP-element group 388:  members (3) 
      -- CP-element group 388: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1171_Update/ack
      -- CP-element group 388: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1171_update_completed_
      -- CP-element group 388: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1171_Update/$exit
      -- 
    ack_2431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 388_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend214_ifx_xthen286_taken_1050_delayed_1_0_1169_inst_ack_1, ack => zeropad3D_CP_676_elements(388)); -- 
    -- CP-element group 389:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	276 
    -- CP-element group 389: 	280 
    -- CP-element group 389: 	284 
    -- CP-element group 389: 	288 
    -- CP-element group 389: 	292 
    -- CP-element group 389: 	296 
    -- CP-element group 389: 	300 
    -- CP-element group 389: 	304 
    -- CP-element group 389: 	308 
    -- CP-element group 389: 	312 
    -- CP-element group 389: 	256 
    -- CP-element group 389: 	264 
    -- CP-element group 389: 	268 
    -- CP-element group 389: marked-predecessors 
    -- CP-element group 389: 	391 
    -- CP-element group 389: successors 
    -- CP-element group 389: 	391 
    -- CP-element group 389:  members (3) 
      -- CP-element group 389: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1179_sample_start_
      -- CP-element group 389: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1179_Sample/$entry
      -- CP-element group 389: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1179_Sample/req
      -- 
    req_2439_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2439_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(389), ack => W_add230_1056_delayed_2_0_1177_inst_req_0); -- 
    zeropad3D_cp_element_group_389: block -- 
      constant place_capacities: IntegerArray(0 to 13) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1);
      constant place_markings: IntegerArray(0 to 13)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 1);
      constant place_delays: IntegerArray(0 to 13) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_389"; 
      signal preds: BooleanArray(1 to 14); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(276) & zeropad3D_CP_676_elements(280) & zeropad3D_CP_676_elements(284) & zeropad3D_CP_676_elements(288) & zeropad3D_CP_676_elements(292) & zeropad3D_CP_676_elements(296) & zeropad3D_CP_676_elements(300) & zeropad3D_CP_676_elements(304) & zeropad3D_CP_676_elements(308) & zeropad3D_CP_676_elements(312) & zeropad3D_CP_676_elements(256) & zeropad3D_CP_676_elements(264) & zeropad3D_CP_676_elements(268) & zeropad3D_CP_676_elements(391);
      gj_zeropad3D_cp_element_group_389 : generic_join generic map(name => joinName, number_of_predecessors => 14, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(389), clk => clk, reset => reset); --
    end block;
    -- CP-element group 390:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: marked-predecessors 
    -- CP-element group 390: 	392 
    -- CP-element group 390: 	395 
    -- CP-element group 390: successors 
    -- CP-element group 390: 	392 
    -- CP-element group 390:  members (3) 
      -- CP-element group 390: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1179_update_start_
      -- CP-element group 390: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1179_Update/$entry
      -- CP-element group 390: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1179_Update/req
      -- 
    req_2444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(390), ack => W_add230_1056_delayed_2_0_1177_inst_req_1); -- 
    zeropad3D_cp_element_group_390: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_390"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(392) & zeropad3D_CP_676_elements(395);
      gj_zeropad3D_cp_element_group_390 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(390), clk => clk, reset => reset); --
    end block;
    -- CP-element group 391:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: 	389 
    -- CP-element group 391: successors 
    -- CP-element group 391: marked-successors 
    -- CP-element group 391: 	278 
    -- CP-element group 391: 	282 
    -- CP-element group 391: 	389 
    -- CP-element group 391: 	286 
    -- CP-element group 391: 	290 
    -- CP-element group 391: 	294 
    -- CP-element group 391: 	298 
    -- CP-element group 391: 	302 
    -- CP-element group 391: 	306 
    -- CP-element group 391: 	310 
    -- CP-element group 391: 	254 
    -- CP-element group 391: 	262 
    -- CP-element group 391: 	266 
    -- CP-element group 391: 	274 
    -- CP-element group 391:  members (3) 
      -- CP-element group 391: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1179_sample_completed_
      -- CP-element group 391: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1179_Sample/$exit
      -- CP-element group 391: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1179_Sample/ack
      -- 
    ack_2440_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 391_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add230_1056_delayed_2_0_1177_inst_ack_0, ack => zeropad3D_CP_676_elements(391)); -- 
    -- CP-element group 392:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 392: predecessors 
    -- CP-element group 392: 	390 
    -- CP-element group 392: successors 
    -- CP-element group 392: 	393 
    -- CP-element group 392: marked-successors 
    -- CP-element group 392: 	390 
    -- CP-element group 392:  members (3) 
      -- CP-element group 392: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1179_update_completed_
      -- CP-element group 392: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1179_Update/$exit
      -- CP-element group 392: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1179_Update/ack
      -- 
    ack_2445_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 392_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add230_1056_delayed_2_0_1177_inst_ack_1, ack => zeropad3D_CP_676_elements(392)); -- 
    -- CP-element group 393:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 393: predecessors 
    -- CP-element group 393: 	356 
    -- CP-element group 393: 	372 
    -- CP-element group 393: 	384 
    -- CP-element group 393: 	388 
    -- CP-element group 393: 	392 
    -- CP-element group 393: marked-predecessors 
    -- CP-element group 393: 	395 
    -- CP-element group 393: successors 
    -- CP-element group 393: 	395 
    -- CP-element group 393:  members (3) 
      -- CP-element group 393: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1184_sample_start_
      -- CP-element group 393: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1184_Sample/$entry
      -- CP-element group 393: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1184_Sample/rr
      -- 
    rr_2453_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2453_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(393), ack => type_cast_1184_inst_req_0); -- 
    zeropad3D_cp_element_group_393: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_393"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(356) & zeropad3D_CP_676_elements(372) & zeropad3D_CP_676_elements(384) & zeropad3D_CP_676_elements(388) & zeropad3D_CP_676_elements(392) & zeropad3D_CP_676_elements(395);
      gj_zeropad3D_cp_element_group_393 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(393), clk => clk, reset => reset); --
    end block;
    -- CP-element group 394:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 394: predecessors 
    -- CP-element group 394: marked-predecessors 
    -- CP-element group 394: 	396 
    -- CP-element group 394: 	407 
    -- CP-element group 394: successors 
    -- CP-element group 394: 	396 
    -- CP-element group 394:  members (3) 
      -- CP-element group 394: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1184_update_start_
      -- CP-element group 394: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1184_Update/$entry
      -- CP-element group 394: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1184_Update/cr
      -- 
    cr_2458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(394), ack => type_cast_1184_inst_req_1); -- 
    zeropad3D_cp_element_group_394: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_394"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(396) & zeropad3D_CP_676_elements(407);
      gj_zeropad3D_cp_element_group_394 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(394), clk => clk, reset => reset); --
    end block;
    -- CP-element group 395:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 395: predecessors 
    -- CP-element group 395: 	393 
    -- CP-element group 395: successors 
    -- CP-element group 395: marked-successors 
    -- CP-element group 395: 	354 
    -- CP-element group 395: 	370 
    -- CP-element group 395: 	382 
    -- CP-element group 395: 	386 
    -- CP-element group 395: 	390 
    -- CP-element group 395: 	393 
    -- CP-element group 395:  members (3) 
      -- CP-element group 395: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1184_sample_completed_
      -- CP-element group 395: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1184_Sample/$exit
      -- CP-element group 395: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1184_Sample/ra
      -- 
    ra_2454_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 395_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1184_inst_ack_0, ack => zeropad3D_CP_676_elements(395)); -- 
    -- CP-element group 396:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 396: predecessors 
    -- CP-element group 396: 	394 
    -- CP-element group 396: successors 
    -- CP-element group 396: 	405 
    -- CP-element group 396: marked-successors 
    -- CP-element group 396: 	394 
    -- CP-element group 396:  members (3) 
      -- CP-element group 396: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1184_update_completed_
      -- CP-element group 396: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1184_Update/$exit
      -- CP-element group 396: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1184_Update/ca
      -- 
    ca_2459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 396_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1184_inst_ack_1, ack => zeropad3D_CP_676_elements(396)); -- 
    -- CP-element group 397:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 397: predecessors 
    -- CP-element group 397: 	356 
    -- CP-element group 397: 	372 
    -- CP-element group 397: 	384 
    -- CP-element group 397: 	388 
    -- CP-element group 397: marked-predecessors 
    -- CP-element group 397: 	399 
    -- CP-element group 397: successors 
    -- CP-element group 397: 	399 
    -- CP-element group 397:  members (3) 
      -- CP-element group 397: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1188_sample_start_
      -- CP-element group 397: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1188_Sample/$entry
      -- CP-element group 397: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1188_Sample/req
      -- 
    req_2467_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2467_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(397), ack => W_ifx_xthen286_exec_guard_1060_delayed_1_0_1186_inst_req_0); -- 
    zeropad3D_cp_element_group_397: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_397"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(356) & zeropad3D_CP_676_elements(372) & zeropad3D_CP_676_elements(384) & zeropad3D_CP_676_elements(388) & zeropad3D_CP_676_elements(399);
      gj_zeropad3D_cp_element_group_397 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(397), clk => clk, reset => reset); --
    end block;
    -- CP-element group 398:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 398: predecessors 
    -- CP-element group 398: marked-predecessors 
    -- CP-element group 398: 	400 
    -- CP-element group 398: successors 
    -- CP-element group 398: 	400 
    -- CP-element group 398:  members (3) 
      -- CP-element group 398: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1188_update_start_
      -- CP-element group 398: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1188_Update/$entry
      -- CP-element group 398: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1188_Update/req
      -- 
    req_2472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(398), ack => W_ifx_xthen286_exec_guard_1060_delayed_1_0_1186_inst_req_1); -- 
    zeropad3D_cp_element_group_398: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_398"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad3D_CP_676_elements(400);
      gj_zeropad3D_cp_element_group_398 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(398), clk => clk, reset => reset); --
    end block;
    -- CP-element group 399:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 399: predecessors 
    -- CP-element group 399: 	397 
    -- CP-element group 399: successors 
    -- CP-element group 399: marked-successors 
    -- CP-element group 399: 	354 
    -- CP-element group 399: 	370 
    -- CP-element group 399: 	382 
    -- CP-element group 399: 	386 
    -- CP-element group 399: 	397 
    -- CP-element group 399:  members (3) 
      -- CP-element group 399: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1188_sample_completed_
      -- CP-element group 399: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1188_Sample/$exit
      -- CP-element group 399: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1188_Sample/ack
      -- 
    ack_2468_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 399_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen286_exec_guard_1060_delayed_1_0_1186_inst_ack_0, ack => zeropad3D_CP_676_elements(399)); -- 
    -- CP-element group 400:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 400: predecessors 
    -- CP-element group 400: 	398 
    -- CP-element group 400: successors 
    -- CP-element group 400: 	496 
    -- CP-element group 400: marked-successors 
    -- CP-element group 400: 	398 
    -- CP-element group 400:  members (3) 
      -- CP-element group 400: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1188_update_completed_
      -- CP-element group 400: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1188_Update/$exit
      -- CP-element group 400: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1188_Update/ack
      -- 
    ack_2473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 400_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen286_exec_guard_1060_delayed_1_0_1186_inst_ack_1, ack => zeropad3D_CP_676_elements(400)); -- 
    -- CP-element group 401:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 401: predecessors 
    -- CP-element group 401: 	356 
    -- CP-element group 401: 	372 
    -- CP-element group 401: 	384 
    -- CP-element group 401: 	388 
    -- CP-element group 401: marked-predecessors 
    -- CP-element group 401: 	403 
    -- CP-element group 401: successors 
    -- CP-element group 401: 	403 
    -- CP-element group 401:  members (3) 
      -- CP-element group 401: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1201_sample_start_
      -- CP-element group 401: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1201_Sample/$entry
      -- CP-element group 401: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1201_Sample/req
      -- 
    req_2481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(401), ack => W_ifx_xthen286_exec_guard_1070_delayed_1_0_1199_inst_req_0); -- 
    zeropad3D_cp_element_group_401: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_401"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(356) & zeropad3D_CP_676_elements(372) & zeropad3D_CP_676_elements(384) & zeropad3D_CP_676_elements(388) & zeropad3D_CP_676_elements(403);
      gj_zeropad3D_cp_element_group_401 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(401), clk => clk, reset => reset); --
    end block;
    -- CP-element group 402:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 402: predecessors 
    -- CP-element group 402: marked-predecessors 
    -- CP-element group 402: 	404 
    -- CP-element group 402: 	407 
    -- CP-element group 402: successors 
    -- CP-element group 402: 	404 
    -- CP-element group 402:  members (3) 
      -- CP-element group 402: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1201_update_start_
      -- CP-element group 402: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1201_Update/$entry
      -- CP-element group 402: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1201_Update/req
      -- 
    req_2486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(402), ack => W_ifx_xthen286_exec_guard_1070_delayed_1_0_1199_inst_req_1); -- 
    zeropad3D_cp_element_group_402: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_402"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(404) & zeropad3D_CP_676_elements(407);
      gj_zeropad3D_cp_element_group_402 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(402), clk => clk, reset => reset); --
    end block;
    -- CP-element group 403:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 403: predecessors 
    -- CP-element group 403: 	401 
    -- CP-element group 403: successors 
    -- CP-element group 403: marked-successors 
    -- CP-element group 403: 	354 
    -- CP-element group 403: 	370 
    -- CP-element group 403: 	382 
    -- CP-element group 403: 	386 
    -- CP-element group 403: 	401 
    -- CP-element group 403:  members (3) 
      -- CP-element group 403: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1201_sample_completed_
      -- CP-element group 403: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1201_Sample/$exit
      -- CP-element group 403: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1201_Sample/ack
      -- 
    ack_2482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 403_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen286_exec_guard_1070_delayed_1_0_1199_inst_ack_0, ack => zeropad3D_CP_676_elements(403)); -- 
    -- CP-element group 404:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 404: predecessors 
    -- CP-element group 404: 	402 
    -- CP-element group 404: successors 
    -- CP-element group 404: 	405 
    -- CP-element group 404: marked-successors 
    -- CP-element group 404: 	402 
    -- CP-element group 404:  members (3) 
      -- CP-element group 404: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1201_update_completed_
      -- CP-element group 404: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1201_Update/$exit
      -- CP-element group 404: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1201_Update/ack
      -- 
    ack_2487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 404_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen286_exec_guard_1070_delayed_1_0_1199_inst_ack_1, ack => zeropad3D_CP_676_elements(404)); -- 
    -- CP-element group 405:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 405: predecessors 
    -- CP-element group 405: 	396 
    -- CP-element group 405: 	404 
    -- CP-element group 405: marked-predecessors 
    -- CP-element group 405: 	407 
    -- CP-element group 405: successors 
    -- CP-element group 405: 	407 
    -- CP-element group 405:  members (3) 
      -- CP-element group 405: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1206_sample_start_
      -- CP-element group 405: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1206_Sample/$entry
      -- CP-element group 405: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1206_Sample/rr
      -- 
    rr_2495_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2495_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(405), ack => type_cast_1206_inst_req_0); -- 
    zeropad3D_cp_element_group_405: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_405"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(396) & zeropad3D_CP_676_elements(404) & zeropad3D_CP_676_elements(407);
      gj_zeropad3D_cp_element_group_405 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(405), clk => clk, reset => reset); --
    end block;
    -- CP-element group 406:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 406: predecessors 
    -- CP-element group 406: marked-predecessors 
    -- CP-element group 406: 	408 
    -- CP-element group 406: 	412 
    -- CP-element group 406: successors 
    -- CP-element group 406: 	408 
    -- CP-element group 406:  members (3) 
      -- CP-element group 406: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1206_update_start_
      -- CP-element group 406: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1206_Update/$entry
      -- CP-element group 406: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1206_Update/cr
      -- 
    cr_2500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(406), ack => type_cast_1206_inst_req_1); -- 
    zeropad3D_cp_element_group_406: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_406"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(408) & zeropad3D_CP_676_elements(412);
      gj_zeropad3D_cp_element_group_406 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(406), clk => clk, reset => reset); --
    end block;
    -- CP-element group 407:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 407: predecessors 
    -- CP-element group 407: 	405 
    -- CP-element group 407: successors 
    -- CP-element group 407: marked-successors 
    -- CP-element group 407: 	394 
    -- CP-element group 407: 	402 
    -- CP-element group 407: 	405 
    -- CP-element group 407:  members (3) 
      -- CP-element group 407: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1206_sample_completed_
      -- CP-element group 407: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1206_Sample/$exit
      -- CP-element group 407: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1206_Sample/ra
      -- 
    ra_2496_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 407_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1206_inst_ack_0, ack => zeropad3D_CP_676_elements(407)); -- 
    -- CP-element group 408:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 408: predecessors 
    -- CP-element group 408: 	406 
    -- CP-element group 408: successors 
    -- CP-element group 408: 	412 
    -- CP-element group 408: marked-successors 
    -- CP-element group 408: 	406 
    -- CP-element group 408:  members (16) 
      -- CP-element group 408: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1206_update_completed_
      -- CP-element group 408: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1206_Update/$exit
      -- CP-element group 408: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1206_Update/ca
      -- CP-element group 408: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1212_index_resized_1
      -- CP-element group 408: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1212_index_scaled_1
      -- CP-element group 408: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1212_index_computed_1
      -- CP-element group 408: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1212_index_resize_1/$entry
      -- CP-element group 408: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1212_index_resize_1/$exit
      -- CP-element group 408: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1212_index_resize_1/index_resize_req
      -- CP-element group 408: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1212_index_resize_1/index_resize_ack
      -- CP-element group 408: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1212_index_scale_1/$entry
      -- CP-element group 408: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1212_index_scale_1/$exit
      -- CP-element group 408: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1212_index_scale_1/scale_rename_req
      -- CP-element group 408: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1212_index_scale_1/scale_rename_ack
      -- CP-element group 408: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1212_final_index_sum_regn_Sample/$entry
      -- CP-element group 408: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1212_final_index_sum_regn_Sample/req
      -- 
    ca_2501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 408_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1206_inst_ack_1, ack => zeropad3D_CP_676_elements(408)); -- 
    req_2526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(408), ack => array_obj_ref_1212_index_offset_req_0); -- 
    -- CP-element group 409:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 409: predecessors 
    -- CP-element group 409: 	413 
    -- CP-element group 409: marked-predecessors 
    -- CP-element group 409: 	414 
    -- CP-element group 409: successors 
    -- CP-element group 409: 	414 
    -- CP-element group 409:  members (3) 
      -- CP-element group 409: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/addr_of_1213_sample_start_
      -- CP-element group 409: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/addr_of_1213_request/$entry
      -- CP-element group 409: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/addr_of_1213_request/req
      -- 
    req_2541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(409), ack => addr_of_1213_final_reg_req_0); -- 
    zeropad3D_cp_element_group_409: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_409"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(413) & zeropad3D_CP_676_elements(414);
      gj_zeropad3D_cp_element_group_409 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(409), clk => clk, reset => reset); --
    end block;
    -- CP-element group 410:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 410: predecessors 
    -- CP-element group 410: 	134 
    -- CP-element group 410: marked-predecessors 
    -- CP-element group 410: 	415 
    -- CP-element group 410: 	418 
    -- CP-element group 410: successors 
    -- CP-element group 410: 	415 
    -- CP-element group 410:  members (3) 
      -- CP-element group 410: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/addr_of_1213_update_start_
      -- CP-element group 410: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/addr_of_1213_complete/$entry
      -- CP-element group 410: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/addr_of_1213_complete/req
      -- 
    req_2546_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2546_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(410), ack => addr_of_1213_final_reg_req_1); -- 
    zeropad3D_cp_element_group_410: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_410"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(134) & zeropad3D_CP_676_elements(415) & zeropad3D_CP_676_elements(418);
      gj_zeropad3D_cp_element_group_410 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(410), clk => clk, reset => reset); --
    end block;
    -- CP-element group 411:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 411: predecessors 
    -- CP-element group 411: 	134 
    -- CP-element group 411: marked-predecessors 
    -- CP-element group 411: 	413 
    -- CP-element group 411: 	414 
    -- CP-element group 411: successors 
    -- CP-element group 411: 	413 
    -- CP-element group 411:  members (3) 
      -- CP-element group 411: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1212_final_index_sum_regn_update_start
      -- CP-element group 411: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1212_final_index_sum_regn_Update/$entry
      -- CP-element group 411: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1212_final_index_sum_regn_Update/req
      -- 
    req_2531_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2531_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(411), ack => array_obj_ref_1212_index_offset_req_1); -- 
    zeropad3D_cp_element_group_411: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_411"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(134) & zeropad3D_CP_676_elements(413) & zeropad3D_CP_676_elements(414);
      gj_zeropad3D_cp_element_group_411 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(411), clk => clk, reset => reset); --
    end block;
    -- CP-element group 412:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 412: predecessors 
    -- CP-element group 412: 	408 
    -- CP-element group 412: successors 
    -- CP-element group 412: 	496 
    -- CP-element group 412: marked-successors 
    -- CP-element group 412: 	406 
    -- CP-element group 412:  members (3) 
      -- CP-element group 412: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1212_final_index_sum_regn_sample_complete
      -- CP-element group 412: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1212_final_index_sum_regn_Sample/$exit
      -- CP-element group 412: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1212_final_index_sum_regn_Sample/ack
      -- 
    ack_2527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 412_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1212_index_offset_ack_0, ack => zeropad3D_CP_676_elements(412)); -- 
    -- CP-element group 413:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 413: predecessors 
    -- CP-element group 413: 	411 
    -- CP-element group 413: successors 
    -- CP-element group 413: 	409 
    -- CP-element group 413: marked-successors 
    -- CP-element group 413: 	411 
    -- CP-element group 413:  members (8) 
      -- CP-element group 413: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1212_root_address_calculated
      -- CP-element group 413: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1212_offset_calculated
      -- CP-element group 413: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1212_final_index_sum_regn_Update/$exit
      -- CP-element group 413: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1212_final_index_sum_regn_Update/ack
      -- CP-element group 413: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1212_base_plus_offset/$entry
      -- CP-element group 413: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1212_base_plus_offset/$exit
      -- CP-element group 413: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1212_base_plus_offset/sum_rename_req
      -- CP-element group 413: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1212_base_plus_offset/sum_rename_ack
      -- 
    ack_2532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 413_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1212_index_offset_ack_1, ack => zeropad3D_CP_676_elements(413)); -- 
    -- CP-element group 414:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 414: predecessors 
    -- CP-element group 414: 	409 
    -- CP-element group 414: successors 
    -- CP-element group 414: marked-successors 
    -- CP-element group 414: 	409 
    -- CP-element group 414: 	411 
    -- CP-element group 414:  members (3) 
      -- CP-element group 414: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/addr_of_1213_sample_completed_
      -- CP-element group 414: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/addr_of_1213_request/$exit
      -- CP-element group 414: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/addr_of_1213_request/ack
      -- 
    ack_2542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 414_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1213_final_reg_ack_0, ack => zeropad3D_CP_676_elements(414)); -- 
    -- CP-element group 415:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 415: predecessors 
    -- CP-element group 415: 	410 
    -- CP-element group 415: successors 
    -- CP-element group 415: 	416 
    -- CP-element group 415: marked-successors 
    -- CP-element group 415: 	410 
    -- CP-element group 415:  members (19) 
      -- CP-element group 415: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/addr_of_1213_update_completed_
      -- CP-element group 415: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/addr_of_1213_complete/$exit
      -- CP-element group 415: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/addr_of_1213_complete/ack
      -- CP-element group 415: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1217_base_address_calculated
      -- CP-element group 415: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1217_word_address_calculated
      -- CP-element group 415: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1217_root_address_calculated
      -- CP-element group 415: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1217_base_address_resized
      -- CP-element group 415: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1217_base_addr_resize/$entry
      -- CP-element group 415: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1217_base_addr_resize/$exit
      -- CP-element group 415: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1217_base_addr_resize/base_resize_req
      -- CP-element group 415: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1217_base_addr_resize/base_resize_ack
      -- CP-element group 415: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1217_base_plus_offset/$entry
      -- CP-element group 415: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1217_base_plus_offset/$exit
      -- CP-element group 415: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1217_base_plus_offset/sum_rename_req
      -- CP-element group 415: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1217_base_plus_offset/sum_rename_ack
      -- CP-element group 415: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1217_word_addrgen/$entry
      -- CP-element group 415: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1217_word_addrgen/$exit
      -- CP-element group 415: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1217_word_addrgen/root_register_req
      -- CP-element group 415: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1217_word_addrgen/root_register_ack
      -- 
    ack_2547_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 415_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1213_final_reg_ack_1, ack => zeropad3D_CP_676_elements(415)); -- 
    -- CP-element group 416:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 416: predecessors 
    -- CP-element group 416: 	415 
    -- CP-element group 416: marked-predecessors 
    -- CP-element group 416: 	418 
    -- CP-element group 416: 	492 
    -- CP-element group 416: successors 
    -- CP-element group 416: 	418 
    -- CP-element group 416:  members (9) 
      -- CP-element group 416: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1217_sample_start_
      -- CP-element group 416: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1217_Sample/$entry
      -- CP-element group 416: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1217_Sample/ptr_deref_1217_Split/$entry
      -- CP-element group 416: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1217_Sample/ptr_deref_1217_Split/$exit
      -- CP-element group 416: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1217_Sample/ptr_deref_1217_Split/split_req
      -- CP-element group 416: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1217_Sample/ptr_deref_1217_Split/split_ack
      -- CP-element group 416: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1217_Sample/word_access_start/$entry
      -- CP-element group 416: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1217_Sample/word_access_start/word_0/$entry
      -- CP-element group 416: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1217_Sample/word_access_start/word_0/rr
      -- 
    rr_2585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(416), ack => ptr_deref_1217_store_0_req_0); -- 
    zeropad3D_cp_element_group_416: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_416"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(415) & zeropad3D_CP_676_elements(418) & zeropad3D_CP_676_elements(492);
      gj_zeropad3D_cp_element_group_416 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(416), clk => clk, reset => reset); --
    end block;
    -- CP-element group 417:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 417: predecessors 
    -- CP-element group 417: marked-predecessors 
    -- CP-element group 417: 	419 
    -- CP-element group 417: successors 
    -- CP-element group 417: 	419 
    -- CP-element group 417:  members (5) 
      -- CP-element group 417: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1217_update_start_
      -- CP-element group 417: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1217_Update/$entry
      -- CP-element group 417: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1217_Update/word_access_complete/$entry
      -- CP-element group 417: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1217_Update/word_access_complete/word_0/$entry
      -- CP-element group 417: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1217_Update/word_access_complete/word_0/cr
      -- 
    cr_2596_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2596_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(417), ack => ptr_deref_1217_store_0_req_1); -- 
    zeropad3D_cp_element_group_417: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_417"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad3D_CP_676_elements(419);
      gj_zeropad3D_cp_element_group_417 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(417), clk => clk, reset => reset); --
    end block;
    -- CP-element group 418:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 418: predecessors 
    -- CP-element group 418: 	416 
    -- CP-element group 418: successors 
    -- CP-element group 418: 	495 
    -- CP-element group 418: marked-successors 
    -- CP-element group 418: 	410 
    -- CP-element group 418: 	416 
    -- CP-element group 418:  members (5) 
      -- CP-element group 418: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1217_sample_completed_
      -- CP-element group 418: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1217_Sample/$exit
      -- CP-element group 418: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1217_Sample/word_access_start/$exit
      -- CP-element group 418: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1217_Sample/word_access_start/word_0/$exit
      -- CP-element group 418: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1217_Sample/word_access_start/word_0/ra
      -- 
    ra_2586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 418_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1217_store_0_ack_0, ack => zeropad3D_CP_676_elements(418)); -- 
    -- CP-element group 419:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 419: predecessors 
    -- CP-element group 419: 	417 
    -- CP-element group 419: successors 
    -- CP-element group 419: 	496 
    -- CP-element group 419: marked-successors 
    -- CP-element group 419: 	417 
    -- CP-element group 419:  members (5) 
      -- CP-element group 419: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1217_update_completed_
      -- CP-element group 419: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1217_Update/$exit
      -- CP-element group 419: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1217_Update/word_access_complete/$exit
      -- CP-element group 419: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1217_Update/word_access_complete/word_0/$exit
      -- CP-element group 419: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1217_Update/word_access_complete/word_0/ca
      -- 
    ca_2597_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 419_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1217_store_0_ack_1, ack => zeropad3D_CP_676_elements(419)); -- 
    -- CP-element group 420:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 420: predecessors 
    -- CP-element group 420: 	276 
    -- CP-element group 420: 	280 
    -- CP-element group 420: 	284 
    -- CP-element group 420: 	288 
    -- CP-element group 420: 	292 
    -- CP-element group 420: 	296 
    -- CP-element group 420: 	300 
    -- CP-element group 420: 	304 
    -- CP-element group 420: 	308 
    -- CP-element group 420: 	312 
    -- CP-element group 420: 	256 
    -- CP-element group 420: 	264 
    -- CP-element group 420: 	268 
    -- CP-element group 420: marked-predecessors 
    -- CP-element group 420: 	422 
    -- CP-element group 420: successors 
    -- CP-element group 420: 	422 
    -- CP-element group 420:  members (3) 
      -- CP-element group 420: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1226_sample_start_
      -- CP-element group 420: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1226_Sample/$entry
      -- CP-element group 420: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1226_Sample/req
      -- 
    req_2605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(420), ack => W_add252_1094_delayed_2_0_1224_inst_req_0); -- 
    zeropad3D_cp_element_group_420: block -- 
      constant place_capacities: IntegerArray(0 to 13) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1);
      constant place_markings: IntegerArray(0 to 13)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 1);
      constant place_delays: IntegerArray(0 to 13) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_420"; 
      signal preds: BooleanArray(1 to 14); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(276) & zeropad3D_CP_676_elements(280) & zeropad3D_CP_676_elements(284) & zeropad3D_CP_676_elements(288) & zeropad3D_CP_676_elements(292) & zeropad3D_CP_676_elements(296) & zeropad3D_CP_676_elements(300) & zeropad3D_CP_676_elements(304) & zeropad3D_CP_676_elements(308) & zeropad3D_CP_676_elements(312) & zeropad3D_CP_676_elements(256) & zeropad3D_CP_676_elements(264) & zeropad3D_CP_676_elements(268) & zeropad3D_CP_676_elements(422);
      gj_zeropad3D_cp_element_group_420 : generic_join generic map(name => joinName, number_of_predecessors => 14, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(420), clk => clk, reset => reset); --
    end block;
    -- CP-element group 421:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 421: predecessors 
    -- CP-element group 421: marked-predecessors 
    -- CP-element group 421: 	423 
    -- CP-element group 421: 	426 
    -- CP-element group 421: successors 
    -- CP-element group 421: 	423 
    -- CP-element group 421:  members (3) 
      -- CP-element group 421: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1226_update_start_
      -- CP-element group 421: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1226_Update/$entry
      -- CP-element group 421: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1226_Update/req
      -- 
    req_2610_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2610_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(421), ack => W_add252_1094_delayed_2_0_1224_inst_req_1); -- 
    zeropad3D_cp_element_group_421: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_421"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(423) & zeropad3D_CP_676_elements(426);
      gj_zeropad3D_cp_element_group_421 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(421), clk => clk, reset => reset); --
    end block;
    -- CP-element group 422:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 422: predecessors 
    -- CP-element group 422: 	420 
    -- CP-element group 422: successors 
    -- CP-element group 422: marked-successors 
    -- CP-element group 422: 	278 
    -- CP-element group 422: 	282 
    -- CP-element group 422: 	286 
    -- CP-element group 422: 	420 
    -- CP-element group 422: 	290 
    -- CP-element group 422: 	294 
    -- CP-element group 422: 	298 
    -- CP-element group 422: 	302 
    -- CP-element group 422: 	306 
    -- CP-element group 422: 	310 
    -- CP-element group 422: 	254 
    -- CP-element group 422: 	262 
    -- CP-element group 422: 	266 
    -- CP-element group 422: 	274 
    -- CP-element group 422:  members (3) 
      -- CP-element group 422: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1226_sample_completed_
      -- CP-element group 422: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1226_Sample/$exit
      -- CP-element group 422: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1226_Sample/ack
      -- 
    ack_2606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 422_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add252_1094_delayed_2_0_1224_inst_ack_0, ack => zeropad3D_CP_676_elements(422)); -- 
    -- CP-element group 423:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 423: predecessors 
    -- CP-element group 423: 	421 
    -- CP-element group 423: successors 
    -- CP-element group 423: 	424 
    -- CP-element group 423: marked-successors 
    -- CP-element group 423: 	421 
    -- CP-element group 423:  members (3) 
      -- CP-element group 423: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1226_update_completed_
      -- CP-element group 423: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1226_Update/$exit
      -- CP-element group 423: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1226_Update/ack
      -- 
    ack_2611_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 423_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add252_1094_delayed_2_0_1224_inst_ack_1, ack => zeropad3D_CP_676_elements(423)); -- 
    -- CP-element group 424:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 424: predecessors 
    -- CP-element group 424: 	356 
    -- CP-element group 424: 	372 
    -- CP-element group 424: 	380 
    -- CP-element group 424: 	423 
    -- CP-element group 424: marked-predecessors 
    -- CP-element group 424: 	426 
    -- CP-element group 424: successors 
    -- CP-element group 424: 	426 
    -- CP-element group 424:  members (3) 
      -- CP-element group 424: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1231_sample_start_
      -- CP-element group 424: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1231_Sample/$entry
      -- CP-element group 424: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1231_Sample/rr
      -- 
    rr_2619_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2619_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(424), ack => type_cast_1231_inst_req_0); -- 
    zeropad3D_cp_element_group_424: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_424"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(356) & zeropad3D_CP_676_elements(372) & zeropad3D_CP_676_elements(380) & zeropad3D_CP_676_elements(423) & zeropad3D_CP_676_elements(426);
      gj_zeropad3D_cp_element_group_424 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(424), clk => clk, reset => reset); --
    end block;
    -- CP-element group 425:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 425: predecessors 
    -- CP-element group 425: marked-predecessors 
    -- CP-element group 425: 	427 
    -- CP-element group 425: 	438 
    -- CP-element group 425: successors 
    -- CP-element group 425: 	427 
    -- CP-element group 425:  members (3) 
      -- CP-element group 425: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1231_update_start_
      -- CP-element group 425: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1231_Update/$entry
      -- CP-element group 425: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1231_Update/cr
      -- 
    cr_2624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(425), ack => type_cast_1231_inst_req_1); -- 
    zeropad3D_cp_element_group_425: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_425"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(427) & zeropad3D_CP_676_elements(438);
      gj_zeropad3D_cp_element_group_425 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(425), clk => clk, reset => reset); --
    end block;
    -- CP-element group 426:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 426: predecessors 
    -- CP-element group 426: 	424 
    -- CP-element group 426: successors 
    -- CP-element group 426: marked-successors 
    -- CP-element group 426: 	354 
    -- CP-element group 426: 	370 
    -- CP-element group 426: 	378 
    -- CP-element group 426: 	421 
    -- CP-element group 426: 	424 
    -- CP-element group 426:  members (3) 
      -- CP-element group 426: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1231_sample_completed_
      -- CP-element group 426: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1231_Sample/$exit
      -- CP-element group 426: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1231_Sample/ra
      -- 
    ra_2620_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 426_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1231_inst_ack_0, ack => zeropad3D_CP_676_elements(426)); -- 
    -- CP-element group 427:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 427: predecessors 
    -- CP-element group 427: 	425 
    -- CP-element group 427: successors 
    -- CP-element group 427: 	436 
    -- CP-element group 427: marked-successors 
    -- CP-element group 427: 	425 
    -- CP-element group 427:  members (3) 
      -- CP-element group 427: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1231_update_completed_
      -- CP-element group 427: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1231_Update/$exit
      -- CP-element group 427: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1231_Update/ca
      -- 
    ca_2625_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 427_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1231_inst_ack_1, ack => zeropad3D_CP_676_elements(427)); -- 
    -- CP-element group 428:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 428: predecessors 
    -- CP-element group 428: 	356 
    -- CP-element group 428: 	372 
    -- CP-element group 428: 	380 
    -- CP-element group 428: marked-predecessors 
    -- CP-element group 428: 	430 
    -- CP-element group 428: successors 
    -- CP-element group 428: 	430 
    -- CP-element group 428:  members (3) 
      -- CP-element group 428: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1235_sample_start_
      -- CP-element group 428: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1235_Sample/$entry
      -- CP-element group 428: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1235_Sample/req
      -- 
    req_2633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(428), ack => W_ifx_xelse292_exec_guard_1098_delayed_1_0_1233_inst_req_0); -- 
    zeropad3D_cp_element_group_428: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_428"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(356) & zeropad3D_CP_676_elements(372) & zeropad3D_CP_676_elements(380) & zeropad3D_CP_676_elements(430);
      gj_zeropad3D_cp_element_group_428 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(428), clk => clk, reset => reset); --
    end block;
    -- CP-element group 429:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 429: predecessors 
    -- CP-element group 429: marked-predecessors 
    -- CP-element group 429: 	431 
    -- CP-element group 429: successors 
    -- CP-element group 429: 	431 
    -- CP-element group 429:  members (3) 
      -- CP-element group 429: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1235_update_start_
      -- CP-element group 429: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1235_Update/$entry
      -- CP-element group 429: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1235_Update/req
      -- 
    req_2638_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2638_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(429), ack => W_ifx_xelse292_exec_guard_1098_delayed_1_0_1233_inst_req_1); -- 
    zeropad3D_cp_element_group_429: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_429"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad3D_CP_676_elements(431);
      gj_zeropad3D_cp_element_group_429 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(429), clk => clk, reset => reset); --
    end block;
    -- CP-element group 430:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 430: predecessors 
    -- CP-element group 430: 	428 
    -- CP-element group 430: successors 
    -- CP-element group 430: marked-successors 
    -- CP-element group 430: 	354 
    -- CP-element group 430: 	370 
    -- CP-element group 430: 	378 
    -- CP-element group 430: 	428 
    -- CP-element group 430:  members (3) 
      -- CP-element group 430: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1235_sample_completed_
      -- CP-element group 430: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1235_Sample/$exit
      -- CP-element group 430: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1235_Sample/ack
      -- 
    ack_2634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 430_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse292_exec_guard_1098_delayed_1_0_1233_inst_ack_0, ack => zeropad3D_CP_676_elements(430)); -- 
    -- CP-element group 431:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 431: predecessors 
    -- CP-element group 431: 	429 
    -- CP-element group 431: successors 
    -- CP-element group 431: 	496 
    -- CP-element group 431: marked-successors 
    -- CP-element group 431: 	429 
    -- CP-element group 431:  members (3) 
      -- CP-element group 431: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1235_update_completed_
      -- CP-element group 431: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1235_Update/$exit
      -- CP-element group 431: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1235_Update/ack
      -- 
    ack_2639_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 431_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse292_exec_guard_1098_delayed_1_0_1233_inst_ack_1, ack => zeropad3D_CP_676_elements(431)); -- 
    -- CP-element group 432:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 432: predecessors 
    -- CP-element group 432: 	356 
    -- CP-element group 432: 	372 
    -- CP-element group 432: 	380 
    -- CP-element group 432: marked-predecessors 
    -- CP-element group 432: 	434 
    -- CP-element group 432: successors 
    -- CP-element group 432: 	434 
    -- CP-element group 432:  members (3) 
      -- CP-element group 432: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1248_sample_start_
      -- CP-element group 432: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1248_Sample/$entry
      -- CP-element group 432: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1248_Sample/req
      -- 
    req_2647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(432), ack => W_ifx_xelse292_exec_guard_1108_delayed_1_0_1246_inst_req_0); -- 
    zeropad3D_cp_element_group_432: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_432"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(356) & zeropad3D_CP_676_elements(372) & zeropad3D_CP_676_elements(380) & zeropad3D_CP_676_elements(434);
      gj_zeropad3D_cp_element_group_432 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(432), clk => clk, reset => reset); --
    end block;
    -- CP-element group 433:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 433: predecessors 
    -- CP-element group 433: marked-predecessors 
    -- CP-element group 433: 	435 
    -- CP-element group 433: 	438 
    -- CP-element group 433: successors 
    -- CP-element group 433: 	435 
    -- CP-element group 433:  members (3) 
      -- CP-element group 433: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1248_update_start_
      -- CP-element group 433: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1248_Update/$entry
      -- CP-element group 433: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1248_Update/req
      -- 
    req_2652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(433), ack => W_ifx_xelse292_exec_guard_1108_delayed_1_0_1246_inst_req_1); -- 
    zeropad3D_cp_element_group_433: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_433"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(435) & zeropad3D_CP_676_elements(438);
      gj_zeropad3D_cp_element_group_433 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(433), clk => clk, reset => reset); --
    end block;
    -- CP-element group 434:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 434: predecessors 
    -- CP-element group 434: 	432 
    -- CP-element group 434: successors 
    -- CP-element group 434: marked-successors 
    -- CP-element group 434: 	354 
    -- CP-element group 434: 	370 
    -- CP-element group 434: 	378 
    -- CP-element group 434: 	432 
    -- CP-element group 434:  members (3) 
      -- CP-element group 434: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1248_sample_completed_
      -- CP-element group 434: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1248_Sample/$exit
      -- CP-element group 434: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1248_Sample/ack
      -- 
    ack_2648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 434_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse292_exec_guard_1108_delayed_1_0_1246_inst_ack_0, ack => zeropad3D_CP_676_elements(434)); -- 
    -- CP-element group 435:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 435: predecessors 
    -- CP-element group 435: 	433 
    -- CP-element group 435: successors 
    -- CP-element group 435: 	436 
    -- CP-element group 435: marked-successors 
    -- CP-element group 435: 	433 
    -- CP-element group 435:  members (3) 
      -- CP-element group 435: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1248_update_completed_
      -- CP-element group 435: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1248_Update/$exit
      -- CP-element group 435: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1248_Update/ack
      -- 
    ack_2653_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 435_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse292_exec_guard_1108_delayed_1_0_1246_inst_ack_1, ack => zeropad3D_CP_676_elements(435)); -- 
    -- CP-element group 436:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 436: predecessors 
    -- CP-element group 436: 	427 
    -- CP-element group 436: 	435 
    -- CP-element group 436: marked-predecessors 
    -- CP-element group 436: 	438 
    -- CP-element group 436: successors 
    -- CP-element group 436: 	438 
    -- CP-element group 436:  members (3) 
      -- CP-element group 436: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1253_sample_start_
      -- CP-element group 436: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1253_Sample/$entry
      -- CP-element group 436: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1253_Sample/rr
      -- 
    rr_2661_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2661_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(436), ack => type_cast_1253_inst_req_0); -- 
    zeropad3D_cp_element_group_436: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_436"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(427) & zeropad3D_CP_676_elements(435) & zeropad3D_CP_676_elements(438);
      gj_zeropad3D_cp_element_group_436 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(436), clk => clk, reset => reset); --
    end block;
    -- CP-element group 437:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 437: predecessors 
    -- CP-element group 437: marked-predecessors 
    -- CP-element group 437: 	439 
    -- CP-element group 437: 	443 
    -- CP-element group 437: successors 
    -- CP-element group 437: 	439 
    -- CP-element group 437:  members (3) 
      -- CP-element group 437: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1253_update_start_
      -- CP-element group 437: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1253_Update/$entry
      -- CP-element group 437: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1253_Update/cr
      -- 
    cr_2666_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2666_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(437), ack => type_cast_1253_inst_req_1); -- 
    zeropad3D_cp_element_group_437: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_437"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(439) & zeropad3D_CP_676_elements(443);
      gj_zeropad3D_cp_element_group_437 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(437), clk => clk, reset => reset); --
    end block;
    -- CP-element group 438:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 438: predecessors 
    -- CP-element group 438: 	436 
    -- CP-element group 438: successors 
    -- CP-element group 438: marked-successors 
    -- CP-element group 438: 	425 
    -- CP-element group 438: 	433 
    -- CP-element group 438: 	436 
    -- CP-element group 438:  members (3) 
      -- CP-element group 438: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1253_sample_completed_
      -- CP-element group 438: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1253_Sample/$exit
      -- CP-element group 438: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1253_Sample/ra
      -- 
    ra_2662_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 438_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1253_inst_ack_0, ack => zeropad3D_CP_676_elements(438)); -- 
    -- CP-element group 439:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 439: predecessors 
    -- CP-element group 439: 	437 
    -- CP-element group 439: successors 
    -- CP-element group 439: 	443 
    -- CP-element group 439: marked-successors 
    -- CP-element group 439: 	437 
    -- CP-element group 439:  members (16) 
      -- CP-element group 439: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1253_update_completed_
      -- CP-element group 439: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1253_Update/$exit
      -- CP-element group 439: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1253_Update/ca
      -- CP-element group 439: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1259_index_resized_1
      -- CP-element group 439: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1259_index_scaled_1
      -- CP-element group 439: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1259_index_computed_1
      -- CP-element group 439: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1259_index_resize_1/$entry
      -- CP-element group 439: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1259_index_resize_1/$exit
      -- CP-element group 439: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1259_index_resize_1/index_resize_req
      -- CP-element group 439: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1259_index_resize_1/index_resize_ack
      -- CP-element group 439: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1259_index_scale_1/$entry
      -- CP-element group 439: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1259_index_scale_1/$exit
      -- CP-element group 439: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1259_index_scale_1/scale_rename_req
      -- CP-element group 439: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1259_index_scale_1/scale_rename_ack
      -- CP-element group 439: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1259_final_index_sum_regn_Sample/$entry
      -- CP-element group 439: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1259_final_index_sum_regn_Sample/req
      -- 
    ca_2667_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 439_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1253_inst_ack_1, ack => zeropad3D_CP_676_elements(439)); -- 
    req_2692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(439), ack => array_obj_ref_1259_index_offset_req_0); -- 
    -- CP-element group 440:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 440: predecessors 
    -- CP-element group 440: 	444 
    -- CP-element group 440: marked-predecessors 
    -- CP-element group 440: 	445 
    -- CP-element group 440: successors 
    -- CP-element group 440: 	445 
    -- CP-element group 440:  members (3) 
      -- CP-element group 440: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/addr_of_1260_sample_start_
      -- CP-element group 440: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/addr_of_1260_request/$entry
      -- CP-element group 440: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/addr_of_1260_request/req
      -- 
    req_2707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(440), ack => addr_of_1260_final_reg_req_0); -- 
    zeropad3D_cp_element_group_440: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_440"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(444) & zeropad3D_CP_676_elements(445);
      gj_zeropad3D_cp_element_group_440 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(440), clk => clk, reset => reset); --
    end block;
    -- CP-element group 441:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 441: predecessors 
    -- CP-element group 441: 	134 
    -- CP-element group 441: marked-predecessors 
    -- CP-element group 441: 	446 
    -- CP-element group 441: 	453 
    -- CP-element group 441: successors 
    -- CP-element group 441: 	446 
    -- CP-element group 441:  members (3) 
      -- CP-element group 441: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/addr_of_1260_update_start_
      -- CP-element group 441: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/addr_of_1260_complete/$entry
      -- CP-element group 441: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/addr_of_1260_complete/req
      -- 
    req_2712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(441), ack => addr_of_1260_final_reg_req_1); -- 
    zeropad3D_cp_element_group_441: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_441"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(134) & zeropad3D_CP_676_elements(446) & zeropad3D_CP_676_elements(453);
      gj_zeropad3D_cp_element_group_441 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(441), clk => clk, reset => reset); --
    end block;
    -- CP-element group 442:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 442: predecessors 
    -- CP-element group 442: 	134 
    -- CP-element group 442: marked-predecessors 
    -- CP-element group 442: 	444 
    -- CP-element group 442: 	445 
    -- CP-element group 442: successors 
    -- CP-element group 442: 	444 
    -- CP-element group 442:  members (3) 
      -- CP-element group 442: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1259_final_index_sum_regn_update_start
      -- CP-element group 442: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1259_final_index_sum_regn_Update/$entry
      -- CP-element group 442: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1259_final_index_sum_regn_Update/req
      -- 
    req_2697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(442), ack => array_obj_ref_1259_index_offset_req_1); -- 
    zeropad3D_cp_element_group_442: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_442"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(134) & zeropad3D_CP_676_elements(444) & zeropad3D_CP_676_elements(445);
      gj_zeropad3D_cp_element_group_442 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(442), clk => clk, reset => reset); --
    end block;
    -- CP-element group 443:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 443: predecessors 
    -- CP-element group 443: 	439 
    -- CP-element group 443: successors 
    -- CP-element group 443: 	496 
    -- CP-element group 443: marked-successors 
    -- CP-element group 443: 	437 
    -- CP-element group 443:  members (3) 
      -- CP-element group 443: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1259_final_index_sum_regn_sample_complete
      -- CP-element group 443: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1259_final_index_sum_regn_Sample/$exit
      -- CP-element group 443: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1259_final_index_sum_regn_Sample/ack
      -- 
    ack_2693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 443_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1259_index_offset_ack_0, ack => zeropad3D_CP_676_elements(443)); -- 
    -- CP-element group 444:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 444: predecessors 
    -- CP-element group 444: 	442 
    -- CP-element group 444: successors 
    -- CP-element group 444: 	440 
    -- CP-element group 444: marked-successors 
    -- CP-element group 444: 	442 
    -- CP-element group 444:  members (8) 
      -- CP-element group 444: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1259_root_address_calculated
      -- CP-element group 444: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1259_offset_calculated
      -- CP-element group 444: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1259_final_index_sum_regn_Update/$exit
      -- CP-element group 444: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1259_final_index_sum_regn_Update/ack
      -- CP-element group 444: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1259_base_plus_offset/$entry
      -- CP-element group 444: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1259_base_plus_offset/$exit
      -- CP-element group 444: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1259_base_plus_offset/sum_rename_req
      -- CP-element group 444: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1259_base_plus_offset/sum_rename_ack
      -- 
    ack_2698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 444_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1259_index_offset_ack_1, ack => zeropad3D_CP_676_elements(444)); -- 
    -- CP-element group 445:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 445: predecessors 
    -- CP-element group 445: 	440 
    -- CP-element group 445: successors 
    -- CP-element group 445: marked-successors 
    -- CP-element group 445: 	440 
    -- CP-element group 445: 	442 
    -- CP-element group 445:  members (3) 
      -- CP-element group 445: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/addr_of_1260_sample_completed_
      -- CP-element group 445: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/addr_of_1260_request/$exit
      -- CP-element group 445: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/addr_of_1260_request/ack
      -- 
    ack_2708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 445_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1260_final_reg_ack_0, ack => zeropad3D_CP_676_elements(445)); -- 
    -- CP-element group 446:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 446: predecessors 
    -- CP-element group 446: 	441 
    -- CP-element group 446: successors 
    -- CP-element group 446: 	451 
    -- CP-element group 446: marked-successors 
    -- CP-element group 446: 	441 
    -- CP-element group 446:  members (19) 
      -- CP-element group 446: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1268_base_plus_offset/sum_rename_req
      -- CP-element group 446: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1268_word_addrgen/root_register_req
      -- CP-element group 446: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1268_word_addrgen/$exit
      -- CP-element group 446: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1268_word_addrgen/$entry
      -- CP-element group 446: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1268_base_addr_resize/$entry
      -- CP-element group 446: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1268_base_addr_resize/$exit
      -- CP-element group 446: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1268_base_address_resized
      -- CP-element group 446: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1268_base_plus_offset/sum_rename_ack
      -- CP-element group 446: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1268_base_addr_resize/base_resize_req
      -- CP-element group 446: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1268_base_plus_offset/$entry
      -- CP-element group 446: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1268_base_addr_resize/base_resize_ack
      -- CP-element group 446: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1268_base_plus_offset/$exit
      -- CP-element group 446: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1268_root_address_calculated
      -- CP-element group 446: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1268_word_address_calculated
      -- CP-element group 446: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1268_base_address_calculated
      -- CP-element group 446: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1268_word_addrgen/root_register_ack
      -- CP-element group 446: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/addr_of_1260_update_completed_
      -- CP-element group 446: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/addr_of_1260_complete/$exit
      -- CP-element group 446: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/addr_of_1260_complete/ack
      -- 
    ack_2713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 446_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1260_final_reg_ack_1, ack => zeropad3D_CP_676_elements(446)); -- 
    -- CP-element group 447:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 447: predecessors 
    -- CP-element group 447: 	356 
    -- CP-element group 447: 	372 
    -- CP-element group 447: 	380 
    -- CP-element group 447: marked-predecessors 
    -- CP-element group 447: 	449 
    -- CP-element group 447: successors 
    -- CP-element group 447: 	449 
    -- CP-element group 447:  members (3) 
      -- CP-element group 447: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1264_sample_start_
      -- CP-element group 447: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1264_Sample/$entry
      -- CP-element group 447: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1264_Sample/req
      -- 
    req_2721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(447), ack => W_ifx_xelse292_exec_guard_1121_delayed_8_0_1262_inst_req_0); -- 
    zeropad3D_cp_element_group_447: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_447"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(356) & zeropad3D_CP_676_elements(372) & zeropad3D_CP_676_elements(380) & zeropad3D_CP_676_elements(449);
      gj_zeropad3D_cp_element_group_447 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(447), clk => clk, reset => reset); --
    end block;
    -- CP-element group 448:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 448: predecessors 
    -- CP-element group 448: marked-predecessors 
    -- CP-element group 448: 	450 
    -- CP-element group 448: 	453 
    -- CP-element group 448: successors 
    -- CP-element group 448: 	450 
    -- CP-element group 448:  members (3) 
      -- CP-element group 448: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1264_update_start_
      -- CP-element group 448: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1264_Update/$entry
      -- CP-element group 448: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1264_Update/req
      -- 
    req_2726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(448), ack => W_ifx_xelse292_exec_guard_1121_delayed_8_0_1262_inst_req_1); -- 
    zeropad3D_cp_element_group_448: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_448"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(450) & zeropad3D_CP_676_elements(453);
      gj_zeropad3D_cp_element_group_448 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(448), clk => clk, reset => reset); --
    end block;
    -- CP-element group 449:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 449: predecessors 
    -- CP-element group 449: 	447 
    -- CP-element group 449: successors 
    -- CP-element group 449: marked-successors 
    -- CP-element group 449: 	354 
    -- CP-element group 449: 	370 
    -- CP-element group 449: 	378 
    -- CP-element group 449: 	447 
    -- CP-element group 449:  members (3) 
      -- CP-element group 449: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1264_sample_completed_
      -- CP-element group 449: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1264_Sample/$exit
      -- CP-element group 449: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1264_Sample/ack
      -- 
    ack_2722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 449_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse292_exec_guard_1121_delayed_8_0_1262_inst_ack_0, ack => zeropad3D_CP_676_elements(449)); -- 
    -- CP-element group 450:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 450: predecessors 
    -- CP-element group 450: 	448 
    -- CP-element group 450: successors 
    -- CP-element group 450: 	451 
    -- CP-element group 450: marked-successors 
    -- CP-element group 450: 	448 
    -- CP-element group 450:  members (3) 
      -- CP-element group 450: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1264_update_completed_
      -- CP-element group 450: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1264_Update/$exit
      -- CP-element group 450: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1264_Update/ack
      -- 
    ack_2727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 450_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse292_exec_guard_1121_delayed_8_0_1262_inst_ack_1, ack => zeropad3D_CP_676_elements(450)); -- 
    -- CP-element group 451:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 451: predecessors 
    -- CP-element group 451: 	446 
    -- CP-element group 451: 	450 
    -- CP-element group 451: marked-predecessors 
    -- CP-element group 451: 	453 
    -- CP-element group 451: successors 
    -- CP-element group 451: 	453 
    -- CP-element group 451:  members (5) 
      -- CP-element group 451: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1268_Sample/word_access_start/$entry
      -- CP-element group 451: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1268_Sample/word_access_start/word_0/rr
      -- CP-element group 451: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1268_Sample/word_access_start/word_0/$entry
      -- CP-element group 451: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1268_Sample/$entry
      -- CP-element group 451: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1268_sample_start_
      -- 
    rr_2760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(451), ack => ptr_deref_1268_load_0_req_0); -- 
    zeropad3D_cp_element_group_451: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_451"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(446) & zeropad3D_CP_676_elements(450) & zeropad3D_CP_676_elements(453);
      gj_zeropad3D_cp_element_group_451 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(451), clk => clk, reset => reset); --
    end block;
    -- CP-element group 452:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 452: predecessors 
    -- CP-element group 452: marked-predecessors 
    -- CP-element group 452: 	454 
    -- CP-element group 452: 	492 
    -- CP-element group 452: successors 
    -- CP-element group 452: 	454 
    -- CP-element group 452:  members (5) 
      -- CP-element group 452: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1268_Update/word_access_complete/word_0/cr
      -- CP-element group 452: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1268_Update/word_access_complete/word_0/$entry
      -- CP-element group 452: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1268_Update/word_access_complete/$entry
      -- CP-element group 452: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1268_Update/$entry
      -- CP-element group 452: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1268_update_start_
      -- 
    cr_2771_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2771_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(452), ack => ptr_deref_1268_load_0_req_1); -- 
    zeropad3D_cp_element_group_452: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_452"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(454) & zeropad3D_CP_676_elements(492);
      gj_zeropad3D_cp_element_group_452 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(452), clk => clk, reset => reset); --
    end block;
    -- CP-element group 453:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 453: predecessors 
    -- CP-element group 453: 	451 
    -- CP-element group 453: successors 
    -- CP-element group 453: marked-successors 
    -- CP-element group 453: 	441 
    -- CP-element group 453: 	448 
    -- CP-element group 453: 	451 
    -- CP-element group 453:  members (5) 
      -- CP-element group 453: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1268_Sample/word_access_start/word_0/ra
      -- CP-element group 453: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1268_Sample/word_access_start/word_0/$exit
      -- CP-element group 453: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1268_Sample/word_access_start/$exit
      -- CP-element group 453: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1268_Sample/$exit
      -- CP-element group 453: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1268_sample_completed_
      -- 
    ra_2761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 453_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1268_load_0_ack_0, ack => zeropad3D_CP_676_elements(453)); -- 
    -- CP-element group 454:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 454: predecessors 
    -- CP-element group 454: 	452 
    -- CP-element group 454: successors 
    -- CP-element group 454: 	490 
    -- CP-element group 454: marked-successors 
    -- CP-element group 454: 	452 
    -- CP-element group 454:  members (9) 
      -- CP-element group 454: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1268_Update/ptr_deref_1268_Merge/merge_ack
      -- CP-element group 454: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1268_Update/ptr_deref_1268_Merge/merge_req
      -- CP-element group 454: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1268_Update/ptr_deref_1268_Merge/$exit
      -- CP-element group 454: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1268_Update/ptr_deref_1268_Merge/$entry
      -- CP-element group 454: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1268_Update/word_access_complete/word_0/ca
      -- CP-element group 454: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1268_Update/word_access_complete/word_0/$exit
      -- CP-element group 454: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1268_Update/word_access_complete/$exit
      -- CP-element group 454: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1268_Update/$exit
      -- CP-element group 454: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1268_update_completed_
      -- 
    ca_2772_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 454_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1268_load_0_ack_1, ack => zeropad3D_CP_676_elements(454)); -- 
    -- CP-element group 455:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 455: predecessors 
    -- CP-element group 455: 	276 
    -- CP-element group 455: 	280 
    -- CP-element group 455: 	284 
    -- CP-element group 455: 	288 
    -- CP-element group 455: 	292 
    -- CP-element group 455: 	296 
    -- CP-element group 455: 	300 
    -- CP-element group 455: 	304 
    -- CP-element group 455: 	308 
    -- CP-element group 455: 	312 
    -- CP-element group 455: 	256 
    -- CP-element group 455: 	264 
    -- CP-element group 455: 	268 
    -- CP-element group 455: marked-predecessors 
    -- CP-element group 455: 	457 
    -- CP-element group 455: successors 
    -- CP-element group 455: 	457 
    -- CP-element group 455:  members (3) 
      -- CP-element group 455: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1272_Sample/$entry
      -- CP-element group 455: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1272_Sample/req
      -- CP-element group 455: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1272_sample_start_
      -- 
    req_2785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(455), ack => W_add230_1128_delayed_2_0_1270_inst_req_0); -- 
    zeropad3D_cp_element_group_455: block -- 
      constant place_capacities: IntegerArray(0 to 13) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1);
      constant place_markings: IntegerArray(0 to 13)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 1);
      constant place_delays: IntegerArray(0 to 13) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_455"; 
      signal preds: BooleanArray(1 to 14); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(276) & zeropad3D_CP_676_elements(280) & zeropad3D_CP_676_elements(284) & zeropad3D_CP_676_elements(288) & zeropad3D_CP_676_elements(292) & zeropad3D_CP_676_elements(296) & zeropad3D_CP_676_elements(300) & zeropad3D_CP_676_elements(304) & zeropad3D_CP_676_elements(308) & zeropad3D_CP_676_elements(312) & zeropad3D_CP_676_elements(256) & zeropad3D_CP_676_elements(264) & zeropad3D_CP_676_elements(268) & zeropad3D_CP_676_elements(457);
      gj_zeropad3D_cp_element_group_455 : generic_join generic map(name => joinName, number_of_predecessors => 14, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(455), clk => clk, reset => reset); --
    end block;
    -- CP-element group 456:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 456: predecessors 
    -- CP-element group 456: marked-predecessors 
    -- CP-element group 456: 	458 
    -- CP-element group 456: 	461 
    -- CP-element group 456: successors 
    -- CP-element group 456: 	458 
    -- CP-element group 456:  members (3) 
      -- CP-element group 456: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1272_update_start_
      -- CP-element group 456: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1272_Update/$entry
      -- CP-element group 456: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1272_Update/req
      -- 
    req_2790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(456), ack => W_add230_1128_delayed_2_0_1270_inst_req_1); -- 
    zeropad3D_cp_element_group_456: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_456"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(458) & zeropad3D_CP_676_elements(461);
      gj_zeropad3D_cp_element_group_456 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(456), clk => clk, reset => reset); --
    end block;
    -- CP-element group 457:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 457: predecessors 
    -- CP-element group 457: 	455 
    -- CP-element group 457: successors 
    -- CP-element group 457: marked-successors 
    -- CP-element group 457: 	278 
    -- CP-element group 457: 	282 
    -- CP-element group 457: 	286 
    -- CP-element group 457: 	290 
    -- CP-element group 457: 	455 
    -- CP-element group 457: 	294 
    -- CP-element group 457: 	298 
    -- CP-element group 457: 	302 
    -- CP-element group 457: 	306 
    -- CP-element group 457: 	310 
    -- CP-element group 457: 	254 
    -- CP-element group 457: 	262 
    -- CP-element group 457: 	266 
    -- CP-element group 457: 	274 
    -- CP-element group 457:  members (3) 
      -- CP-element group 457: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1272_Sample/$exit
      -- CP-element group 457: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1272_Sample/ack
      -- CP-element group 457: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1272_sample_completed_
      -- 
    ack_2786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 457_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add230_1128_delayed_2_0_1270_inst_ack_0, ack => zeropad3D_CP_676_elements(457)); -- 
    -- CP-element group 458:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 458: predecessors 
    -- CP-element group 458: 	456 
    -- CP-element group 458: successors 
    -- CP-element group 458: 	459 
    -- CP-element group 458: marked-successors 
    -- CP-element group 458: 	456 
    -- CP-element group 458:  members (3) 
      -- CP-element group 458: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1272_Update/ack
      -- CP-element group 458: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1272_update_completed_
      -- CP-element group 458: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1272_Update/$exit
      -- 
    ack_2791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 458_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add230_1128_delayed_2_0_1270_inst_ack_1, ack => zeropad3D_CP_676_elements(458)); -- 
    -- CP-element group 459:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 459: predecessors 
    -- CP-element group 459: 	356 
    -- CP-element group 459: 	372 
    -- CP-element group 459: 	380 
    -- CP-element group 459: 	458 
    -- CP-element group 459: marked-predecessors 
    -- CP-element group 459: 	461 
    -- CP-element group 459: successors 
    -- CP-element group 459: 	461 
    -- CP-element group 459:  members (3) 
      -- CP-element group 459: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1277_sample_start_
      -- CP-element group 459: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1277_Sample/$entry
      -- CP-element group 459: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1277_Sample/rr
      -- 
    rr_2799_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2799_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(459), ack => type_cast_1277_inst_req_0); -- 
    zeropad3D_cp_element_group_459: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_459"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(356) & zeropad3D_CP_676_elements(372) & zeropad3D_CP_676_elements(380) & zeropad3D_CP_676_elements(458) & zeropad3D_CP_676_elements(461);
      gj_zeropad3D_cp_element_group_459 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(459), clk => clk, reset => reset); --
    end block;
    -- CP-element group 460:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 460: predecessors 
    -- CP-element group 460: marked-predecessors 
    -- CP-element group 460: 	462 
    -- CP-element group 460: 	473 
    -- CP-element group 460: successors 
    -- CP-element group 460: 	462 
    -- CP-element group 460:  members (3) 
      -- CP-element group 460: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1277_Update/$entry
      -- CP-element group 460: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1277_Update/cr
      -- CP-element group 460: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1277_update_start_
      -- 
    cr_2804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(460), ack => type_cast_1277_inst_req_1); -- 
    zeropad3D_cp_element_group_460: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_460"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(462) & zeropad3D_CP_676_elements(473);
      gj_zeropad3D_cp_element_group_460 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(460), clk => clk, reset => reset); --
    end block;
    -- CP-element group 461:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 461: predecessors 
    -- CP-element group 461: 	459 
    -- CP-element group 461: successors 
    -- CP-element group 461: marked-successors 
    -- CP-element group 461: 	354 
    -- CP-element group 461: 	370 
    -- CP-element group 461: 	378 
    -- CP-element group 461: 	456 
    -- CP-element group 461: 	459 
    -- CP-element group 461:  members (3) 
      -- CP-element group 461: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1277_sample_completed_
      -- CP-element group 461: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1277_Sample/ra
      -- CP-element group 461: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1277_Sample/$exit
      -- 
    ra_2800_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 461_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1277_inst_ack_0, ack => zeropad3D_CP_676_elements(461)); -- 
    -- CP-element group 462:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 462: predecessors 
    -- CP-element group 462: 	460 
    -- CP-element group 462: successors 
    -- CP-element group 462: 	471 
    -- CP-element group 462: marked-successors 
    -- CP-element group 462: 	460 
    -- CP-element group 462:  members (3) 
      -- CP-element group 462: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1277_Update/ca
      -- CP-element group 462: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1277_Update/$exit
      -- CP-element group 462: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1277_update_completed_
      -- 
    ca_2805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 462_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1277_inst_ack_1, ack => zeropad3D_CP_676_elements(462)); -- 
    -- CP-element group 463:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 463: predecessors 
    -- CP-element group 463: 	356 
    -- CP-element group 463: 	372 
    -- CP-element group 463: 	380 
    -- CP-element group 463: marked-predecessors 
    -- CP-element group 463: 	465 
    -- CP-element group 463: successors 
    -- CP-element group 463: 	465 
    -- CP-element group 463:  members (3) 
      -- CP-element group 463: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1281_sample_start_
      -- CP-element group 463: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1281_Sample/req
      -- CP-element group 463: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1281_Sample/$entry
      -- 
    req_2813_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2813_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(463), ack => W_ifx_xelse292_exec_guard_1132_delayed_1_0_1279_inst_req_0); -- 
    zeropad3D_cp_element_group_463: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_463"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(356) & zeropad3D_CP_676_elements(372) & zeropad3D_CP_676_elements(380) & zeropad3D_CP_676_elements(465);
      gj_zeropad3D_cp_element_group_463 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(463), clk => clk, reset => reset); --
    end block;
    -- CP-element group 464:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 464: predecessors 
    -- CP-element group 464: marked-predecessors 
    -- CP-element group 464: 	466 
    -- CP-element group 464: successors 
    -- CP-element group 464: 	466 
    -- CP-element group 464:  members (3) 
      -- CP-element group 464: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1281_Update/req
      -- CP-element group 464: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1281_Update/$entry
      -- CP-element group 464: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1281_update_start_
      -- 
    req_2818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(464), ack => W_ifx_xelse292_exec_guard_1132_delayed_1_0_1279_inst_req_1); -- 
    zeropad3D_cp_element_group_464: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_464"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad3D_CP_676_elements(466);
      gj_zeropad3D_cp_element_group_464 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(464), clk => clk, reset => reset); --
    end block;
    -- CP-element group 465:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 465: predecessors 
    -- CP-element group 465: 	463 
    -- CP-element group 465: successors 
    -- CP-element group 465: marked-successors 
    -- CP-element group 465: 	354 
    -- CP-element group 465: 	370 
    -- CP-element group 465: 	378 
    -- CP-element group 465: 	463 
    -- CP-element group 465:  members (3) 
      -- CP-element group 465: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1281_sample_completed_
      -- CP-element group 465: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1281_Sample/ack
      -- CP-element group 465: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1281_Sample/$exit
      -- 
    ack_2814_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 465_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse292_exec_guard_1132_delayed_1_0_1279_inst_ack_0, ack => zeropad3D_CP_676_elements(465)); -- 
    -- CP-element group 466:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 466: predecessors 
    -- CP-element group 466: 	464 
    -- CP-element group 466: successors 
    -- CP-element group 466: 	496 
    -- CP-element group 466: marked-successors 
    -- CP-element group 466: 	464 
    -- CP-element group 466:  members (3) 
      -- CP-element group 466: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1281_Update/ack
      -- CP-element group 466: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1281_Update/$exit
      -- CP-element group 466: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1281_update_completed_
      -- 
    ack_2819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 466_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse292_exec_guard_1132_delayed_1_0_1279_inst_ack_1, ack => zeropad3D_CP_676_elements(466)); -- 
    -- CP-element group 467:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 467: predecessors 
    -- CP-element group 467: 	356 
    -- CP-element group 467: 	372 
    -- CP-element group 467: 	380 
    -- CP-element group 467: marked-predecessors 
    -- CP-element group 467: 	469 
    -- CP-element group 467: successors 
    -- CP-element group 467: 	469 
    -- CP-element group 467:  members (3) 
      -- CP-element group 467: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1294_Sample/req
      -- CP-element group 467: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1294_Sample/$entry
      -- CP-element group 467: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1294_sample_start_
      -- 
    req_2827_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2827_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(467), ack => W_ifx_xelse292_exec_guard_1142_delayed_1_0_1292_inst_req_0); -- 
    zeropad3D_cp_element_group_467: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_467"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(356) & zeropad3D_CP_676_elements(372) & zeropad3D_CP_676_elements(380) & zeropad3D_CP_676_elements(469);
      gj_zeropad3D_cp_element_group_467 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(467), clk => clk, reset => reset); --
    end block;
    -- CP-element group 468:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 468: predecessors 
    -- CP-element group 468: marked-predecessors 
    -- CP-element group 468: 	470 
    -- CP-element group 468: 	473 
    -- CP-element group 468: successors 
    -- CP-element group 468: 	470 
    -- CP-element group 468:  members (3) 
      -- CP-element group 468: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1294_Update/$entry
      -- CP-element group 468: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1294_Update/req
      -- CP-element group 468: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1294_update_start_
      -- 
    req_2832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(468), ack => W_ifx_xelse292_exec_guard_1142_delayed_1_0_1292_inst_req_1); -- 
    zeropad3D_cp_element_group_468: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_468"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(470) & zeropad3D_CP_676_elements(473);
      gj_zeropad3D_cp_element_group_468 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(468), clk => clk, reset => reset); --
    end block;
    -- CP-element group 469:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 469: predecessors 
    -- CP-element group 469: 	467 
    -- CP-element group 469: successors 
    -- CP-element group 469: marked-successors 
    -- CP-element group 469: 	354 
    -- CP-element group 469: 	370 
    -- CP-element group 469: 	378 
    -- CP-element group 469: 	467 
    -- CP-element group 469:  members (3) 
      -- CP-element group 469: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1294_Sample/ack
      -- CP-element group 469: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1294_Sample/$exit
      -- CP-element group 469: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1294_sample_completed_
      -- 
    ack_2828_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 469_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse292_exec_guard_1142_delayed_1_0_1292_inst_ack_0, ack => zeropad3D_CP_676_elements(469)); -- 
    -- CP-element group 470:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 470: predecessors 
    -- CP-element group 470: 	468 
    -- CP-element group 470: successors 
    -- CP-element group 470: 	471 
    -- CP-element group 470: marked-successors 
    -- CP-element group 470: 	468 
    -- CP-element group 470:  members (3) 
      -- CP-element group 470: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1294_Update/$exit
      -- CP-element group 470: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1294_Update/ack
      -- CP-element group 470: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1294_update_completed_
      -- 
    ack_2833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 470_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse292_exec_guard_1142_delayed_1_0_1292_inst_ack_1, ack => zeropad3D_CP_676_elements(470)); -- 
    -- CP-element group 471:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 471: predecessors 
    -- CP-element group 471: 	462 
    -- CP-element group 471: 	470 
    -- CP-element group 471: marked-predecessors 
    -- CP-element group 471: 	473 
    -- CP-element group 471: successors 
    -- CP-element group 471: 	473 
    -- CP-element group 471:  members (3) 
      -- CP-element group 471: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1299_Sample/$entry
      -- CP-element group 471: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1299_Sample/rr
      -- CP-element group 471: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1299_sample_start_
      -- 
    rr_2841_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2841_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(471), ack => type_cast_1299_inst_req_0); -- 
    zeropad3D_cp_element_group_471: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_471"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(462) & zeropad3D_CP_676_elements(470) & zeropad3D_CP_676_elements(473);
      gj_zeropad3D_cp_element_group_471 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(471), clk => clk, reset => reset); --
    end block;
    -- CP-element group 472:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 472: predecessors 
    -- CP-element group 472: marked-predecessors 
    -- CP-element group 472: 	474 
    -- CP-element group 472: 	478 
    -- CP-element group 472: successors 
    -- CP-element group 472: 	474 
    -- CP-element group 472:  members (3) 
      -- CP-element group 472: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1299_Update/cr
      -- CP-element group 472: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1299_update_start_
      -- CP-element group 472: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1299_Update/$entry
      -- 
    cr_2846_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2846_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(472), ack => type_cast_1299_inst_req_1); -- 
    zeropad3D_cp_element_group_472: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_472"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(474) & zeropad3D_CP_676_elements(478);
      gj_zeropad3D_cp_element_group_472 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(472), clk => clk, reset => reset); --
    end block;
    -- CP-element group 473:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 473: predecessors 
    -- CP-element group 473: 	471 
    -- CP-element group 473: successors 
    -- CP-element group 473: marked-successors 
    -- CP-element group 473: 	460 
    -- CP-element group 473: 	468 
    -- CP-element group 473: 	471 
    -- CP-element group 473:  members (3) 
      -- CP-element group 473: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1299_Sample/$exit
      -- CP-element group 473: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1299_sample_completed_
      -- CP-element group 473: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1299_Sample/ra
      -- 
    ra_2842_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 473_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1299_inst_ack_0, ack => zeropad3D_CP_676_elements(473)); -- 
    -- CP-element group 474:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 474: predecessors 
    -- CP-element group 474: 	472 
    -- CP-element group 474: successors 
    -- CP-element group 474: 	478 
    -- CP-element group 474: marked-successors 
    -- CP-element group 474: 	472 
    -- CP-element group 474:  members (16) 
      -- CP-element group 474: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1299_Update/ca
      -- CP-element group 474: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1299_Update/$exit
      -- CP-element group 474: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1305_final_index_sum_regn_Sample/req
      -- CP-element group 474: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/type_cast_1299_update_completed_
      -- CP-element group 474: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1305_index_scale_1/$exit
      -- CP-element group 474: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1305_final_index_sum_regn_Sample/$entry
      -- CP-element group 474: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1305_index_scale_1/scale_rename_req
      -- CP-element group 474: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1305_index_scale_1/scale_rename_ack
      -- CP-element group 474: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1305_index_resized_1
      -- CP-element group 474: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1305_index_scaled_1
      -- CP-element group 474: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1305_index_scale_1/$entry
      -- CP-element group 474: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1305_index_resize_1/index_resize_ack
      -- CP-element group 474: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1305_index_resize_1/index_resize_req
      -- CP-element group 474: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1305_index_resize_1/$exit
      -- CP-element group 474: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1305_index_resize_1/$entry
      -- CP-element group 474: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1305_index_computed_1
      -- 
    ca_2847_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 474_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1299_inst_ack_1, ack => zeropad3D_CP_676_elements(474)); -- 
    req_2872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(474), ack => array_obj_ref_1305_index_offset_req_0); -- 
    -- CP-element group 475:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 475: predecessors 
    -- CP-element group 475: 	479 
    -- CP-element group 475: marked-predecessors 
    -- CP-element group 475: 	480 
    -- CP-element group 475: successors 
    -- CP-element group 475: 	480 
    -- CP-element group 475:  members (3) 
      -- CP-element group 475: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/addr_of_1306_sample_start_
      -- CP-element group 475: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/addr_of_1306_request/req
      -- CP-element group 475: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/addr_of_1306_request/$entry
      -- 
    req_2887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(475), ack => addr_of_1306_final_reg_req_0); -- 
    zeropad3D_cp_element_group_475: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_475"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(479) & zeropad3D_CP_676_elements(480);
      gj_zeropad3D_cp_element_group_475 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(475), clk => clk, reset => reset); --
    end block;
    -- CP-element group 476:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 476: predecessors 
    -- CP-element group 476: 	134 
    -- CP-element group 476: marked-predecessors 
    -- CP-element group 476: 	481 
    -- CP-element group 476: 	488 
    -- CP-element group 476: successors 
    -- CP-element group 476: 	481 
    -- CP-element group 476:  members (3) 
      -- CP-element group 476: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/addr_of_1306_update_start_
      -- CP-element group 476: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/addr_of_1306_complete/req
      -- CP-element group 476: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/addr_of_1306_complete/$entry
      -- 
    req_2892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(476), ack => addr_of_1306_final_reg_req_1); -- 
    zeropad3D_cp_element_group_476: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_476"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(134) & zeropad3D_CP_676_elements(481) & zeropad3D_CP_676_elements(488);
      gj_zeropad3D_cp_element_group_476 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(476), clk => clk, reset => reset); --
    end block;
    -- CP-element group 477:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 477: predecessors 
    -- CP-element group 477: 	134 
    -- CP-element group 477: marked-predecessors 
    -- CP-element group 477: 	479 
    -- CP-element group 477: 	480 
    -- CP-element group 477: successors 
    -- CP-element group 477: 	479 
    -- CP-element group 477:  members (3) 
      -- CP-element group 477: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1305_final_index_sum_regn_update_start
      -- CP-element group 477: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1305_final_index_sum_regn_Update/req
      -- CP-element group 477: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1305_final_index_sum_regn_Update/$entry
      -- 
    req_2877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(477), ack => array_obj_ref_1305_index_offset_req_1); -- 
    zeropad3D_cp_element_group_477: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_477"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(134) & zeropad3D_CP_676_elements(479) & zeropad3D_CP_676_elements(480);
      gj_zeropad3D_cp_element_group_477 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(477), clk => clk, reset => reset); --
    end block;
    -- CP-element group 478:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 478: predecessors 
    -- CP-element group 478: 	474 
    -- CP-element group 478: successors 
    -- CP-element group 478: 	496 
    -- CP-element group 478: marked-successors 
    -- CP-element group 478: 	472 
    -- CP-element group 478:  members (3) 
      -- CP-element group 478: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1305_final_index_sum_regn_Sample/ack
      -- CP-element group 478: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1305_final_index_sum_regn_sample_complete
      -- CP-element group 478: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1305_final_index_sum_regn_Sample/$exit
      -- 
    ack_2873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 478_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1305_index_offset_ack_0, ack => zeropad3D_CP_676_elements(478)); -- 
    -- CP-element group 479:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 479: predecessors 
    -- CP-element group 479: 	477 
    -- CP-element group 479: successors 
    -- CP-element group 479: 	475 
    -- CP-element group 479: marked-successors 
    -- CP-element group 479: 	477 
    -- CP-element group 479:  members (8) 
      -- CP-element group 479: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1305_root_address_calculated
      -- CP-element group 479: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1305_offset_calculated
      -- CP-element group 479: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1305_base_plus_offset/sum_rename_ack
      -- CP-element group 479: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1305_base_plus_offset/sum_rename_req
      -- CP-element group 479: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1305_base_plus_offset/$exit
      -- CP-element group 479: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1305_base_plus_offset/$entry
      -- CP-element group 479: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1305_final_index_sum_regn_Update/ack
      -- CP-element group 479: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/array_obj_ref_1305_final_index_sum_regn_Update/$exit
      -- 
    ack_2878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 479_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1305_index_offset_ack_1, ack => zeropad3D_CP_676_elements(479)); -- 
    -- CP-element group 480:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 480: predecessors 
    -- CP-element group 480: 	475 
    -- CP-element group 480: successors 
    -- CP-element group 480: marked-successors 
    -- CP-element group 480: 	475 
    -- CP-element group 480: 	477 
    -- CP-element group 480:  members (3) 
      -- CP-element group 480: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/addr_of_1306_sample_completed_
      -- CP-element group 480: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/addr_of_1306_request/ack
      -- CP-element group 480: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/addr_of_1306_request/$exit
      -- 
    ack_2888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 480_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1306_final_reg_ack_0, ack => zeropad3D_CP_676_elements(480)); -- 
    -- CP-element group 481:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 481: predecessors 
    -- CP-element group 481: 	476 
    -- CP-element group 481: successors 
    -- CP-element group 481: 	486 
    -- CP-element group 481: marked-successors 
    -- CP-element group 481: 	476 
    -- CP-element group 481:  members (3) 
      -- CP-element group 481: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/addr_of_1306_update_completed_
      -- CP-element group 481: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/addr_of_1306_complete/ack
      -- CP-element group 481: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/addr_of_1306_complete/$exit
      -- 
    ack_2893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 481_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1306_final_reg_ack_1, ack => zeropad3D_CP_676_elements(481)); -- 
    -- CP-element group 482:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 482: predecessors 
    -- CP-element group 482: 	356 
    -- CP-element group 482: 	372 
    -- CP-element group 482: 	380 
    -- CP-element group 482: marked-predecessors 
    -- CP-element group 482: 	484 
    -- CP-element group 482: successors 
    -- CP-element group 482: 	484 
    -- CP-element group 482:  members (3) 
      -- CP-element group 482: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1310_Sample/req
      -- CP-element group 482: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1310_Sample/$entry
      -- CP-element group 482: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1310_sample_start_
      -- 
    req_2901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(482), ack => W_ifx_xelse292_exec_guard_1155_delayed_14_0_1308_inst_req_0); -- 
    zeropad3D_cp_element_group_482: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_482"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(356) & zeropad3D_CP_676_elements(372) & zeropad3D_CP_676_elements(380) & zeropad3D_CP_676_elements(484);
      gj_zeropad3D_cp_element_group_482 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(482), clk => clk, reset => reset); --
    end block;
    -- CP-element group 483:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 483: predecessors 
    -- CP-element group 483: marked-predecessors 
    -- CP-element group 483: 	485 
    -- CP-element group 483: successors 
    -- CP-element group 483: 	485 
    -- CP-element group 483:  members (3) 
      -- CP-element group 483: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1310_Update/req
      -- CP-element group 483: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1310_Update/$entry
      -- CP-element group 483: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1310_update_start_
      -- 
    req_2906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(483), ack => W_ifx_xelse292_exec_guard_1155_delayed_14_0_1308_inst_req_1); -- 
    zeropad3D_cp_element_group_483: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_483"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad3D_CP_676_elements(485);
      gj_zeropad3D_cp_element_group_483 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(483), clk => clk, reset => reset); --
    end block;
    -- CP-element group 484:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 484: predecessors 
    -- CP-element group 484: 	482 
    -- CP-element group 484: successors 
    -- CP-element group 484: marked-successors 
    -- CP-element group 484: 	354 
    -- CP-element group 484: 	370 
    -- CP-element group 484: 	378 
    -- CP-element group 484: 	482 
    -- CP-element group 484:  members (3) 
      -- CP-element group 484: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1310_Sample/ack
      -- CP-element group 484: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1310_Sample/$exit
      -- CP-element group 484: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1310_sample_completed_
      -- 
    ack_2902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 484_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse292_exec_guard_1155_delayed_14_0_1308_inst_ack_0, ack => zeropad3D_CP_676_elements(484)); -- 
    -- CP-element group 485:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 485: predecessors 
    -- CP-element group 485: 	483 
    -- CP-element group 485: successors 
    -- CP-element group 485: 	496 
    -- CP-element group 485: marked-successors 
    -- CP-element group 485: 	483 
    -- CP-element group 485:  members (3) 
      -- CP-element group 485: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1310_Update/ack
      -- CP-element group 485: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1310_Update/$exit
      -- CP-element group 485: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1310_update_completed_
      -- 
    ack_2907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 485_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse292_exec_guard_1155_delayed_14_0_1308_inst_ack_1, ack => zeropad3D_CP_676_elements(485)); -- 
    -- CP-element group 486:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 486: predecessors 
    -- CP-element group 486: 	481 
    -- CP-element group 486: marked-predecessors 
    -- CP-element group 486: 	488 
    -- CP-element group 486: successors 
    -- CP-element group 486: 	488 
    -- CP-element group 486:  members (3) 
      -- CP-element group 486: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1313_Sample/req
      -- CP-element group 486: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1313_Sample/$entry
      -- CP-element group 486: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1313_sample_start_
      -- 
    req_2915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(486), ack => W_arrayidx303_1156_delayed_5_0_1311_inst_req_0); -- 
    zeropad3D_cp_element_group_486: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_486"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(481) & zeropad3D_CP_676_elements(488);
      gj_zeropad3D_cp_element_group_486 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(486), clk => clk, reset => reset); --
    end block;
    -- CP-element group 487:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 487: predecessors 
    -- CP-element group 487: marked-predecessors 
    -- CP-element group 487: 	489 
    -- CP-element group 487: 	492 
    -- CP-element group 487: successors 
    -- CP-element group 487: 	489 
    -- CP-element group 487:  members (3) 
      -- CP-element group 487: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1313_Update/$entry
      -- CP-element group 487: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1313_Update/req
      -- CP-element group 487: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1313_update_start_
      -- 
    req_2920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(487), ack => W_arrayidx303_1156_delayed_5_0_1311_inst_req_1); -- 
    zeropad3D_cp_element_group_487: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_487"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(489) & zeropad3D_CP_676_elements(492);
      gj_zeropad3D_cp_element_group_487 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(487), clk => clk, reset => reset); --
    end block;
    -- CP-element group 488:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 488: predecessors 
    -- CP-element group 488: 	486 
    -- CP-element group 488: successors 
    -- CP-element group 488: marked-successors 
    -- CP-element group 488: 	476 
    -- CP-element group 488: 	486 
    -- CP-element group 488:  members (3) 
      -- CP-element group 488: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1313_Sample/$exit
      -- CP-element group 488: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1313_Sample/ack
      -- CP-element group 488: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1313_sample_completed_
      -- 
    ack_2916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 488_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_arrayidx303_1156_delayed_5_0_1311_inst_ack_0, ack => zeropad3D_CP_676_elements(488)); -- 
    -- CP-element group 489:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 489: predecessors 
    -- CP-element group 489: 	487 
    -- CP-element group 489: successors 
    -- CP-element group 489: 	490 
    -- CP-element group 489: marked-successors 
    -- CP-element group 489: 	487 
    -- CP-element group 489:  members (19) 
      -- CP-element group 489: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1313_update_completed_
      -- CP-element group 489: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1316_word_address_calculated
      -- CP-element group 489: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1313_Update/$exit
      -- CP-element group 489: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1316_root_address_calculated
      -- CP-element group 489: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/assign_stmt_1313_Update/ack
      -- CP-element group 489: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1316_base_address_resized
      -- CP-element group 489: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1316_base_address_calculated
      -- CP-element group 489: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1316_word_addrgen/root_register_ack
      -- CP-element group 489: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1316_word_addrgen/root_register_req
      -- CP-element group 489: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1316_word_addrgen/$exit
      -- CP-element group 489: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1316_word_addrgen/$entry
      -- CP-element group 489: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1316_base_plus_offset/sum_rename_ack
      -- CP-element group 489: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1316_base_plus_offset/sum_rename_req
      -- CP-element group 489: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1316_base_plus_offset/$exit
      -- CP-element group 489: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1316_base_plus_offset/$entry
      -- CP-element group 489: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1316_base_addr_resize/base_resize_ack
      -- CP-element group 489: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1316_base_addr_resize/base_resize_req
      -- CP-element group 489: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1316_base_addr_resize/$exit
      -- CP-element group 489: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1316_base_addr_resize/$entry
      -- 
    ack_2921_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 489_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_arrayidx303_1156_delayed_5_0_1311_inst_ack_1, ack => zeropad3D_CP_676_elements(489)); -- 
    -- CP-element group 490:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 490: predecessors 
    -- CP-element group 490: 	454 
    -- CP-element group 490: 	489 
    -- CP-element group 490: 	495 
    -- CP-element group 490: marked-predecessors 
    -- CP-element group 490: 	492 
    -- CP-element group 490: successors 
    -- CP-element group 490: 	492 
    -- CP-element group 490:  members (9) 
      -- CP-element group 490: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1316_sample_start_
      -- CP-element group 490: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1316_Sample/word_access_start/word_0/rr
      -- CP-element group 490: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1316_Sample/word_access_start/word_0/$entry
      -- CP-element group 490: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1316_Sample/word_access_start/$entry
      -- CP-element group 490: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1316_Sample/ptr_deref_1316_Split/split_ack
      -- CP-element group 490: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1316_Sample/ptr_deref_1316_Split/split_req
      -- CP-element group 490: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1316_Sample/ptr_deref_1316_Split/$exit
      -- CP-element group 490: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1316_Sample/ptr_deref_1316_Split/$entry
      -- CP-element group 490: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1316_Sample/$entry
      -- 
    rr_2959_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2959_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(490), ack => ptr_deref_1316_store_0_req_0); -- 
    zeropad3D_cp_element_group_490: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_490"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(454) & zeropad3D_CP_676_elements(489) & zeropad3D_CP_676_elements(495) & zeropad3D_CP_676_elements(492);
      gj_zeropad3D_cp_element_group_490 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(490), clk => clk, reset => reset); --
    end block;
    -- CP-element group 491:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 491: predecessors 
    -- CP-element group 491: marked-predecessors 
    -- CP-element group 491: 	493 
    -- CP-element group 491: successors 
    -- CP-element group 491: 	493 
    -- CP-element group 491:  members (5) 
      -- CP-element group 491: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1316_Update/word_access_complete/word_0/cr
      -- CP-element group 491: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1316_update_start_
      -- CP-element group 491: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1316_Update/word_access_complete/word_0/$entry
      -- CP-element group 491: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1316_Update/word_access_complete/$entry
      -- CP-element group 491: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1316_Update/$entry
      -- 
    cr_2970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(491), ack => ptr_deref_1316_store_0_req_1); -- 
    zeropad3D_cp_element_group_491: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_491"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad3D_CP_676_elements(493);
      gj_zeropad3D_cp_element_group_491 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(491), clk => clk, reset => reset); --
    end block;
    -- CP-element group 492:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 492: predecessors 
    -- CP-element group 492: 	490 
    -- CP-element group 492: successors 
    -- CP-element group 492: 	496 
    -- CP-element group 492: marked-successors 
    -- CP-element group 492: 	416 
    -- CP-element group 492: 	452 
    -- CP-element group 492: 	487 
    -- CP-element group 492: 	490 
    -- CP-element group 492:  members (6) 
      -- CP-element group 492: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ring_reenable_memory_space_0
      -- CP-element group 492: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1316_sample_completed_
      -- CP-element group 492: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1316_Sample/word_access_start/word_0/ra
      -- CP-element group 492: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1316_Sample/word_access_start/word_0/$exit
      -- CP-element group 492: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1316_Sample/word_access_start/$exit
      -- CP-element group 492: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1316_Sample/$exit
      -- 
    ra_2960_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 492_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1316_store_0_ack_0, ack => zeropad3D_CP_676_elements(492)); -- 
    -- CP-element group 493:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 493: predecessors 
    -- CP-element group 493: 	491 
    -- CP-element group 493: successors 
    -- CP-element group 493: 	496 
    -- CP-element group 493: marked-successors 
    -- CP-element group 493: 	491 
    -- CP-element group 493:  members (5) 
      -- CP-element group 493: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1316_update_completed_
      -- CP-element group 493: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1316_Update/word_access_complete/word_0/ca
      -- CP-element group 493: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1316_Update/word_access_complete/$exit
      -- CP-element group 493: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1316_Update/word_access_complete/word_0/$exit
      -- CP-element group 493: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1316_Update/$exit
      -- 
    ca_2971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 493_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1316_store_0_ack_1, ack => zeropad3D_CP_676_elements(493)); -- 
    -- CP-element group 494:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 494: predecessors 
    -- CP-element group 494: 	134 
    -- CP-element group 494: successors 
    -- CP-element group 494: 	135 
    -- CP-element group 494:  members (1) 
      -- CP-element group 494: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group zeropad3D_CP_676_elements(494) is a control-delay.
    cp_element_494_delay: control_delay_element  generic map(name => " 494_delay", delay_value => 1)  port map(req => zeropad3D_CP_676_elements(134), ack => zeropad3D_CP_676_elements(494), clk => clk, reset =>reset);
    -- CP-element group 495:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 495: predecessors 
    -- CP-element group 495: 	418 
    -- CP-element group 495: successors 
    -- CP-element group 495: 	490 
    -- CP-element group 495:  members (1) 
      -- CP-element group 495: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/ptr_deref_1217_ptr_deref_1316_delay
      -- 
    -- Element group zeropad3D_CP_676_elements(495) is a control-delay.
    cp_element_495_delay: control_delay_element  generic map(name => " 495_delay", delay_value => 1)  port map(req => zeropad3D_CP_676_elements(418), ack => zeropad3D_CP_676_elements(495), clk => clk, reset =>reset);
    -- CP-element group 496:  join  transition  bypass  pipeline-parent 
    -- CP-element group 496: predecessors 
    -- CP-element group 496: 	324 
    -- CP-element group 496: 	328 
    -- CP-element group 496: 	332 
    -- CP-element group 496: 	340 
    -- CP-element group 496: 	360 
    -- CP-element group 496: 	364 
    -- CP-element group 496: 	368 
    -- CP-element group 496: 	376 
    -- CP-element group 496: 	400 
    -- CP-element group 496: 	412 
    -- CP-element group 496: 	419 
    -- CP-element group 496: 	431 
    -- CP-element group 496: 	443 
    -- CP-element group 496: 	466 
    -- CP-element group 496: 	478 
    -- CP-element group 496: 	485 
    -- CP-element group 496: 	492 
    -- CP-element group 496: 	493 
    -- CP-element group 496: 	224 
    -- CP-element group 496: 	236 
    -- CP-element group 496: 	244 
    -- CP-element group 496: 	260 
    -- CP-element group 496: successors 
    -- CP-element group 496: 	131 
    -- CP-element group 496:  members (1) 
      -- CP-element group 496: 	 branch_block_stmt_222/do_while_stmt_707/do_while_stmt_707_loop_body/$exit
      -- 
    zeropad3D_cp_element_group_496: block -- 
      constant place_capacities: IntegerArray(0 to 21) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 15,11 => 15,12 => 15,13 => 15,14 => 15,15 => 15,16 => 15,17 => 15,18 => 15,19 => 15,20 => 15,21 => 15);
      constant place_markings: IntegerArray(0 to 21)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0);
      constant place_delays: IntegerArray(0 to 21) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_496"; 
      signal preds: BooleanArray(1 to 22); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(324) & zeropad3D_CP_676_elements(328) & zeropad3D_CP_676_elements(332) & zeropad3D_CP_676_elements(340) & zeropad3D_CP_676_elements(360) & zeropad3D_CP_676_elements(364) & zeropad3D_CP_676_elements(368) & zeropad3D_CP_676_elements(376) & zeropad3D_CP_676_elements(400) & zeropad3D_CP_676_elements(412) & zeropad3D_CP_676_elements(419) & zeropad3D_CP_676_elements(431) & zeropad3D_CP_676_elements(443) & zeropad3D_CP_676_elements(466) & zeropad3D_CP_676_elements(478) & zeropad3D_CP_676_elements(485) & zeropad3D_CP_676_elements(492) & zeropad3D_CP_676_elements(493) & zeropad3D_CP_676_elements(224) & zeropad3D_CP_676_elements(236) & zeropad3D_CP_676_elements(244) & zeropad3D_CP_676_elements(260);
      gj_zeropad3D_cp_element_group_496 : generic_join generic map(name => joinName, number_of_predecessors => 22, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(496), clk => clk, reset => reset); --
    end block;
    -- CP-element group 497:  transition  input  bypass  pipeline-parent 
    -- CP-element group 497: predecessors 
    -- CP-element group 497: 	130 
    -- CP-element group 497: successors 
    -- CP-element group 497:  members (2) 
      -- CP-element group 497: 	 branch_block_stmt_222/do_while_stmt_707/loop_exit/ack
      -- CP-element group 497: 	 branch_block_stmt_222/do_while_stmt_707/loop_exit/$exit
      -- 
    ack_2978_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 497_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_707_branch_ack_0, ack => zeropad3D_CP_676_elements(497)); -- 
    -- CP-element group 498:  transition  input  bypass  pipeline-parent 
    -- CP-element group 498: predecessors 
    -- CP-element group 498: 	130 
    -- CP-element group 498: successors 
    -- CP-element group 498:  members (2) 
      -- CP-element group 498: 	 branch_block_stmt_222/do_while_stmt_707/loop_taken/ack
      -- CP-element group 498: 	 branch_block_stmt_222/do_while_stmt_707/loop_taken/$exit
      -- 
    ack_2982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 498_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_707_branch_ack_1, ack => zeropad3D_CP_676_elements(498)); -- 
    -- CP-element group 499:  transition  bypass  pipeline-parent 
    -- CP-element group 499: predecessors 
    -- CP-element group 499: 	128 
    -- CP-element group 499: successors 
    -- CP-element group 499: 	1 
    -- CP-element group 499:  members (1) 
      -- CP-element group 499: 	 branch_block_stmt_222/do_while_stmt_707/$exit
      -- 
    zeropad3D_CP_676_elements(499) <= zeropad3D_CP_676_elements(128);
    -- CP-element group 500:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 500: predecessors 
    -- CP-element group 500: 	1 
    -- CP-element group 500: successors 
    -- CP-element group 500: 	502 
    -- CP-element group 500: 	503 
    -- CP-element group 500:  members (18) 
      -- CP-element group 500: 	 branch_block_stmt_222/assign_stmt_1340__entry__
      -- CP-element group 500: 	 branch_block_stmt_222/merge_stmt_1335__exit__
      -- CP-element group 500: 	 branch_block_stmt_222/assign_stmt_1340/type_cast_1339_Sample/$entry
      -- CP-element group 500: 	 branch_block_stmt_222/if_stmt_1331_if_link/$exit
      -- CP-element group 500: 	 branch_block_stmt_222/ifx_xend304_whilex_xend
      -- CP-element group 500: 	 branch_block_stmt_222/if_stmt_1331_if_link/if_choice_transition
      -- CP-element group 500: 	 branch_block_stmt_222/assign_stmt_1340/type_cast_1339_update_start_
      -- CP-element group 500: 	 branch_block_stmt_222/assign_stmt_1340/$entry
      -- CP-element group 500: 	 branch_block_stmt_222/assign_stmt_1340/type_cast_1339_sample_start_
      -- CP-element group 500: 	 branch_block_stmt_222/assign_stmt_1340/type_cast_1339_Update/cr
      -- CP-element group 500: 	 branch_block_stmt_222/assign_stmt_1340/type_cast_1339_Update/$entry
      -- CP-element group 500: 	 branch_block_stmt_222/assign_stmt_1340/type_cast_1339_Sample/rr
      -- CP-element group 500: 	 branch_block_stmt_222/ifx_xend304_whilex_xend_PhiReq/$entry
      -- CP-element group 500: 	 branch_block_stmt_222/ifx_xend304_whilex_xend_PhiReq/$exit
      -- CP-element group 500: 	 branch_block_stmt_222/merge_stmt_1335_PhiReqMerge
      -- CP-element group 500: 	 branch_block_stmt_222/merge_stmt_1335_PhiAck/$entry
      -- CP-element group 500: 	 branch_block_stmt_222/merge_stmt_1335_PhiAck/$exit
      -- CP-element group 500: 	 branch_block_stmt_222/merge_stmt_1335_PhiAck/dummy
      -- 
    if_choice_transition_2996_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 500_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1331_branch_ack_1, ack => zeropad3D_CP_676_elements(500)); -- 
    cr_3017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(500), ack => type_cast_1339_inst_req_1); -- 
    rr_3012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(500), ack => type_cast_1339_inst_req_0); -- 
    -- CP-element group 501:  merge  transition  place  input  bypass 
    -- CP-element group 501: predecessors 
    -- CP-element group 501: 	1 
    -- CP-element group 501: successors 
    -- CP-element group 501:  members (5) 
      -- CP-element group 501: 	 branch_block_stmt_222/merge_stmt_1335__entry__
      -- CP-element group 501: 	 branch_block_stmt_222/if_stmt_1331__exit__
      -- CP-element group 501: 	 branch_block_stmt_222/if_stmt_1331_else_link/$exit
      -- CP-element group 501: 	 branch_block_stmt_222/if_stmt_1331_else_link/else_choice_transition
      -- CP-element group 501: 	 branch_block_stmt_222/merge_stmt_1335_dead_link/$entry
      -- 
    else_choice_transition_3000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 501_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1331_branch_ack_0, ack => zeropad3D_CP_676_elements(501)); -- 
    -- CP-element group 502:  transition  input  bypass 
    -- CP-element group 502: predecessors 
    -- CP-element group 502: 	500 
    -- CP-element group 502: successors 
    -- CP-element group 502:  members (3) 
      -- CP-element group 502: 	 branch_block_stmt_222/assign_stmt_1340/type_cast_1339_Sample/$exit
      -- CP-element group 502: 	 branch_block_stmt_222/assign_stmt_1340/type_cast_1339_sample_completed_
      -- CP-element group 502: 	 branch_block_stmt_222/assign_stmt_1340/type_cast_1339_Sample/ra
      -- 
    ra_3013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 502_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1339_inst_ack_0, ack => zeropad3D_CP_676_elements(502)); -- 
    -- CP-element group 503:  fork  transition  place  input  output  bypass 
    -- CP-element group 503: predecessors 
    -- CP-element group 503: 	500 
    -- CP-element group 503: successors 
    -- CP-element group 503: 	511 
    -- CP-element group 503: 	513 
    -- CP-element group 503: 	519 
    -- CP-element group 503: 	521 
    -- CP-element group 503: 	523 
    -- CP-element group 503: 	515 
    -- CP-element group 503: 	517 
    -- CP-element group 503: 	507 
    -- CP-element group 503: 	509 
    -- CP-element group 503: 	504 
    -- CP-element group 503: 	505 
    -- CP-element group 503:  members (40) 
      -- CP-element group 503: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451__entry__
      -- CP-element group 503: 	 branch_block_stmt_222/assign_stmt_1340__exit__
      -- CP-element group 503: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1376_update_start_
      -- CP-element group 503: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1347_Update/cr
      -- CP-element group 503: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/call_stmt_1343_sample_start_
      -- CP-element group 503: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1347_Update/$entry
      -- CP-element group 503: 	 branch_block_stmt_222/assign_stmt_1340/type_cast_1339_update_completed_
      -- CP-element group 503: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1356_Update/$entry
      -- CP-element group 503: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1386_Update/cr
      -- CP-element group 503: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1347_update_start_
      -- CP-element group 503: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1386_Update/$entry
      -- CP-element group 503: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/$entry
      -- CP-element group 503: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1396_Update/cr
      -- CP-element group 503: 	 branch_block_stmt_222/assign_stmt_1340/$exit
      -- CP-element group 503: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/call_stmt_1343_Update/ccr
      -- CP-element group 503: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1356_update_start_
      -- CP-element group 503: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1396_Update/$entry
      -- CP-element group 503: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1366_Update/cr
      -- CP-element group 503: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1376_Update/cr
      -- CP-element group 503: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1366_Update/$entry
      -- CP-element group 503: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/call_stmt_1343_Update/$entry
      -- CP-element group 503: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1386_update_start_
      -- CP-element group 503: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/call_stmt_1343_Sample/crr
      -- CP-element group 503: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1376_Update/$entry
      -- CP-element group 503: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/call_stmt_1343_Sample/$entry
      -- CP-element group 503: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1366_update_start_
      -- CP-element group 503: 	 branch_block_stmt_222/assign_stmt_1340/type_cast_1339_Update/ca
      -- CP-element group 503: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/call_stmt_1343_update_start_
      -- CP-element group 503: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1396_update_start_
      -- CP-element group 503: 	 branch_block_stmt_222/assign_stmt_1340/type_cast_1339_Update/$exit
      -- CP-element group 503: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1356_Update/cr
      -- CP-element group 503: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1406_update_start_
      -- CP-element group 503: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1406_Update/$entry
      -- CP-element group 503: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1406_Update/cr
      -- CP-element group 503: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1416_update_start_
      -- CP-element group 503: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1416_Update/$entry
      -- CP-element group 503: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1416_Update/cr
      -- CP-element group 503: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1426_update_start_
      -- CP-element group 503: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1426_Update/$entry
      -- CP-element group 503: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1426_Update/cr
      -- 
    ca_3018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 503_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1339_inst_ack_1, ack => zeropad3D_CP_676_elements(503)); -- 
    cr_3048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(503), ack => type_cast_1347_inst_req_1); -- 
    cr_3104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(503), ack => type_cast_1386_inst_req_1); -- 
    cr_3118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(503), ack => type_cast_1396_inst_req_1); -- 
    ccr_3034_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3034_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(503), ack => call_stmt_1343_call_req_1); -- 
    cr_3076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(503), ack => type_cast_1366_inst_req_1); -- 
    cr_3090_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3090_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(503), ack => type_cast_1376_inst_req_1); -- 
    crr_3029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(503), ack => call_stmt_1343_call_req_0); -- 
    cr_3062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(503), ack => type_cast_1356_inst_req_1); -- 
    cr_3132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(503), ack => type_cast_1406_inst_req_1); -- 
    cr_3146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(503), ack => type_cast_1416_inst_req_1); -- 
    cr_3160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(503), ack => type_cast_1426_inst_req_1); -- 
    -- CP-element group 504:  transition  input  bypass 
    -- CP-element group 504: predecessors 
    -- CP-element group 504: 	503 
    -- CP-element group 504: successors 
    -- CP-element group 504:  members (3) 
      -- CP-element group 504: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/call_stmt_1343_sample_completed_
      -- CP-element group 504: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/call_stmt_1343_Sample/cra
      -- CP-element group 504: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/call_stmt_1343_Sample/$exit
      -- 
    cra_3030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 504_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1343_call_ack_0, ack => zeropad3D_CP_676_elements(504)); -- 
    -- CP-element group 505:  transition  input  output  bypass 
    -- CP-element group 505: predecessors 
    -- CP-element group 505: 	503 
    -- CP-element group 505: successors 
    -- CP-element group 505: 	506 
    -- CP-element group 505:  members (6) 
      -- CP-element group 505: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1347_sample_start_
      -- CP-element group 505: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1347_Sample/rr
      -- CP-element group 505: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/call_stmt_1343_Update/cca
      -- CP-element group 505: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/call_stmt_1343_Update/$exit
      -- CP-element group 505: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1347_Sample/$entry
      -- CP-element group 505: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/call_stmt_1343_update_completed_
      -- 
    cca_3035_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 505_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1343_call_ack_1, ack => zeropad3D_CP_676_elements(505)); -- 
    rr_3043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(505), ack => type_cast_1347_inst_req_0); -- 
    -- CP-element group 506:  transition  input  bypass 
    -- CP-element group 506: predecessors 
    -- CP-element group 506: 	505 
    -- CP-element group 506: successors 
    -- CP-element group 506:  members (3) 
      -- CP-element group 506: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1347_sample_completed_
      -- CP-element group 506: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1347_Sample/ra
      -- CP-element group 506: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1347_Sample/$exit
      -- 
    ra_3044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 506_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1347_inst_ack_0, ack => zeropad3D_CP_676_elements(506)); -- 
    -- CP-element group 507:  fork  transition  input  output  bypass 
    -- CP-element group 507: predecessors 
    -- CP-element group 507: 	503 
    -- CP-element group 507: successors 
    -- CP-element group 507: 	510 
    -- CP-element group 507: 	512 
    -- CP-element group 507: 	520 
    -- CP-element group 507: 	522 
    -- CP-element group 507: 	514 
    -- CP-element group 507: 	516 
    -- CP-element group 507: 	518 
    -- CP-element group 507: 	508 
    -- CP-element group 507:  members (27) 
      -- CP-element group 507: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1347_Update/$exit
      -- CP-element group 507: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1356_Sample/$entry
      -- CP-element group 507: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1366_Sample/rr
      -- CP-element group 507: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1356_Sample/rr
      -- CP-element group 507: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1386_sample_start_
      -- CP-element group 507: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1347_update_completed_
      -- CP-element group 507: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1386_Sample/rr
      -- CP-element group 507: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1386_Sample/$entry
      -- CP-element group 507: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1347_Update/ca
      -- CP-element group 507: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1376_sample_start_
      -- CP-element group 507: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1396_Sample/rr
      -- CP-element group 507: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1366_Sample/$entry
      -- CP-element group 507: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1396_sample_start_
      -- CP-element group 507: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1376_Sample/rr
      -- CP-element group 507: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1356_sample_start_
      -- CP-element group 507: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1376_Sample/$entry
      -- CP-element group 507: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1366_sample_start_
      -- CP-element group 507: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1396_Sample/$entry
      -- CP-element group 507: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1406_sample_start_
      -- CP-element group 507: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1406_Sample/$entry
      -- CP-element group 507: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1406_Sample/rr
      -- CP-element group 507: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1416_sample_start_
      -- CP-element group 507: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1416_Sample/$entry
      -- CP-element group 507: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1416_Sample/rr
      -- CP-element group 507: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1426_sample_start_
      -- CP-element group 507: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1426_Sample/$entry
      -- CP-element group 507: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1426_Sample/rr
      -- 
    ca_3049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 507_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1347_inst_ack_1, ack => zeropad3D_CP_676_elements(507)); -- 
    rr_3071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(507), ack => type_cast_1366_inst_req_0); -- 
    rr_3085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(507), ack => type_cast_1376_inst_req_0); -- 
    rr_3099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(507), ack => type_cast_1386_inst_req_0); -- 
    rr_3141_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3141_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(507), ack => type_cast_1416_inst_req_0); -- 
    rr_3155_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3155_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(507), ack => type_cast_1426_inst_req_0); -- 
    rr_3113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(507), ack => type_cast_1396_inst_req_0); -- 
    rr_3127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(507), ack => type_cast_1406_inst_req_0); -- 
    rr_3057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(507), ack => type_cast_1356_inst_req_0); -- 
    -- CP-element group 508:  transition  input  bypass 
    -- CP-element group 508: predecessors 
    -- CP-element group 508: 	507 
    -- CP-element group 508: successors 
    -- CP-element group 508:  members (3) 
      -- CP-element group 508: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1356_Sample/$exit
      -- CP-element group 508: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1356_Sample/ra
      -- CP-element group 508: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1356_sample_completed_
      -- 
    ra_3058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 508_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1356_inst_ack_0, ack => zeropad3D_CP_676_elements(508)); -- 
    -- CP-element group 509:  transition  input  bypass 
    -- CP-element group 509: predecessors 
    -- CP-element group 509: 	503 
    -- CP-element group 509: successors 
    -- CP-element group 509: 	544 
    -- CP-element group 509:  members (3) 
      -- CP-element group 509: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1356_update_completed_
      -- CP-element group 509: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1356_Update/ca
      -- CP-element group 509: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1356_Update/$exit
      -- 
    ca_3063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 509_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1356_inst_ack_1, ack => zeropad3D_CP_676_elements(509)); -- 
    -- CP-element group 510:  transition  input  bypass 
    -- CP-element group 510: predecessors 
    -- CP-element group 510: 	507 
    -- CP-element group 510: successors 
    -- CP-element group 510:  members (3) 
      -- CP-element group 510: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1366_Sample/ra
      -- CP-element group 510: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1366_Sample/$exit
      -- CP-element group 510: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1366_sample_completed_
      -- 
    ra_3072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 510_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1366_inst_ack_0, ack => zeropad3D_CP_676_elements(510)); -- 
    -- CP-element group 511:  transition  input  bypass 
    -- CP-element group 511: predecessors 
    -- CP-element group 511: 	503 
    -- CP-element group 511: successors 
    -- CP-element group 511: 	541 
    -- CP-element group 511:  members (3) 
      -- CP-element group 511: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1366_Update/ca
      -- CP-element group 511: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1366_Update/$exit
      -- CP-element group 511: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1366_update_completed_
      -- 
    ca_3077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 511_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1366_inst_ack_1, ack => zeropad3D_CP_676_elements(511)); -- 
    -- CP-element group 512:  transition  input  bypass 
    -- CP-element group 512: predecessors 
    -- CP-element group 512: 	507 
    -- CP-element group 512: successors 
    -- CP-element group 512:  members (3) 
      -- CP-element group 512: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1376_sample_completed_
      -- CP-element group 512: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1376_Sample/$exit
      -- CP-element group 512: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1376_Sample/ra
      -- 
    ra_3086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 512_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1376_inst_ack_0, ack => zeropad3D_CP_676_elements(512)); -- 
    -- CP-element group 513:  transition  input  bypass 
    -- CP-element group 513: predecessors 
    -- CP-element group 513: 	503 
    -- CP-element group 513: successors 
    -- CP-element group 513: 	538 
    -- CP-element group 513:  members (3) 
      -- CP-element group 513: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1376_Update/ca
      -- CP-element group 513: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1376_Update/$exit
      -- CP-element group 513: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1376_update_completed_
      -- 
    ca_3091_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 513_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1376_inst_ack_1, ack => zeropad3D_CP_676_elements(513)); -- 
    -- CP-element group 514:  transition  input  bypass 
    -- CP-element group 514: predecessors 
    -- CP-element group 514: 	507 
    -- CP-element group 514: successors 
    -- CP-element group 514:  members (3) 
      -- CP-element group 514: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1386_Sample/$exit
      -- CP-element group 514: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1386_Sample/ra
      -- CP-element group 514: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1386_sample_completed_
      -- 
    ra_3100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 514_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1386_inst_ack_0, ack => zeropad3D_CP_676_elements(514)); -- 
    -- CP-element group 515:  transition  input  bypass 
    -- CP-element group 515: predecessors 
    -- CP-element group 515: 	503 
    -- CP-element group 515: successors 
    -- CP-element group 515: 	535 
    -- CP-element group 515:  members (3) 
      -- CP-element group 515: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1386_Update/$exit
      -- CP-element group 515: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1386_update_completed_
      -- CP-element group 515: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1386_Update/ca
      -- 
    ca_3105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 515_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1386_inst_ack_1, ack => zeropad3D_CP_676_elements(515)); -- 
    -- CP-element group 516:  transition  input  bypass 
    -- CP-element group 516: predecessors 
    -- CP-element group 516: 	507 
    -- CP-element group 516: successors 
    -- CP-element group 516:  members (3) 
      -- CP-element group 516: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1396_Sample/ra
      -- CP-element group 516: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1396_sample_completed_
      -- CP-element group 516: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1396_Sample/$exit
      -- 
    ra_3114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 516_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1396_inst_ack_0, ack => zeropad3D_CP_676_elements(516)); -- 
    -- CP-element group 517:  transition  input  bypass 
    -- CP-element group 517: predecessors 
    -- CP-element group 517: 	503 
    -- CP-element group 517: successors 
    -- CP-element group 517: 	532 
    -- CP-element group 517:  members (3) 
      -- CP-element group 517: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1396_Update/ca
      -- CP-element group 517: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1396_update_completed_
      -- CP-element group 517: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1396_Update/$exit
      -- 
    ca_3119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 517_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1396_inst_ack_1, ack => zeropad3D_CP_676_elements(517)); -- 
    -- CP-element group 518:  transition  input  bypass 
    -- CP-element group 518: predecessors 
    -- CP-element group 518: 	507 
    -- CP-element group 518: successors 
    -- CP-element group 518:  members (3) 
      -- CP-element group 518: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1406_sample_completed_
      -- CP-element group 518: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1406_Sample/$exit
      -- CP-element group 518: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1406_Sample/ra
      -- 
    ra_3128_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 518_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1406_inst_ack_0, ack => zeropad3D_CP_676_elements(518)); -- 
    -- CP-element group 519:  transition  input  bypass 
    -- CP-element group 519: predecessors 
    -- CP-element group 519: 	503 
    -- CP-element group 519: successors 
    -- CP-element group 519: 	529 
    -- CP-element group 519:  members (3) 
      -- CP-element group 519: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1406_update_completed_
      -- CP-element group 519: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1406_Update/$exit
      -- CP-element group 519: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1406_Update/ca
      -- 
    ca_3133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 519_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1406_inst_ack_1, ack => zeropad3D_CP_676_elements(519)); -- 
    -- CP-element group 520:  transition  input  bypass 
    -- CP-element group 520: predecessors 
    -- CP-element group 520: 	507 
    -- CP-element group 520: successors 
    -- CP-element group 520:  members (3) 
      -- CP-element group 520: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1416_sample_completed_
      -- CP-element group 520: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1416_Sample/$exit
      -- CP-element group 520: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1416_Sample/ra
      -- 
    ra_3142_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 520_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1416_inst_ack_0, ack => zeropad3D_CP_676_elements(520)); -- 
    -- CP-element group 521:  transition  input  bypass 
    -- CP-element group 521: predecessors 
    -- CP-element group 521: 	503 
    -- CP-element group 521: successors 
    -- CP-element group 521: 	526 
    -- CP-element group 521:  members (3) 
      -- CP-element group 521: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1416_update_completed_
      -- CP-element group 521: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1416_Update/$exit
      -- CP-element group 521: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1416_Update/ca
      -- 
    ca_3147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 521_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1416_inst_ack_1, ack => zeropad3D_CP_676_elements(521)); -- 
    -- CP-element group 522:  transition  input  bypass 
    -- CP-element group 522: predecessors 
    -- CP-element group 522: 	507 
    -- CP-element group 522: successors 
    -- CP-element group 522:  members (3) 
      -- CP-element group 522: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1426_sample_completed_
      -- CP-element group 522: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1426_Sample/$exit
      -- CP-element group 522: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1426_Sample/ra
      -- 
    ra_3156_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 522_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1426_inst_ack_0, ack => zeropad3D_CP_676_elements(522)); -- 
    -- CP-element group 523:  transition  input  output  bypass 
    -- CP-element group 523: predecessors 
    -- CP-element group 523: 	503 
    -- CP-element group 523: successors 
    -- CP-element group 523: 	524 
    -- CP-element group 523:  members (6) 
      -- CP-element group 523: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1426_update_completed_
      -- CP-element group 523: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1426_Update/$exit
      -- CP-element group 523: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/type_cast_1426_Update/ca
      -- CP-element group 523: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1428_sample_start_
      -- CP-element group 523: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1428_Sample/$entry
      -- CP-element group 523: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1428_Sample/req
      -- 
    ca_3161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 523_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1426_inst_ack_1, ack => zeropad3D_CP_676_elements(523)); -- 
    req_3169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(523), ack => WPIPE_zeropad_output_pipe_1428_inst_req_0); -- 
    -- CP-element group 524:  transition  input  output  bypass 
    -- CP-element group 524: predecessors 
    -- CP-element group 524: 	523 
    -- CP-element group 524: successors 
    -- CP-element group 524: 	525 
    -- CP-element group 524:  members (6) 
      -- CP-element group 524: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1428_sample_completed_
      -- CP-element group 524: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1428_update_start_
      -- CP-element group 524: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1428_Sample/$exit
      -- CP-element group 524: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1428_Sample/ack
      -- CP-element group 524: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1428_Update/$entry
      -- CP-element group 524: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1428_Update/req
      -- 
    ack_3170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 524_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_1428_inst_ack_0, ack => zeropad3D_CP_676_elements(524)); -- 
    req_3174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(524), ack => WPIPE_zeropad_output_pipe_1428_inst_req_1); -- 
    -- CP-element group 525:  transition  input  bypass 
    -- CP-element group 525: predecessors 
    -- CP-element group 525: 	524 
    -- CP-element group 525: successors 
    -- CP-element group 525: 	526 
    -- CP-element group 525:  members (3) 
      -- CP-element group 525: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1428_update_completed_
      -- CP-element group 525: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1428_Update/$exit
      -- CP-element group 525: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1428_Update/ack
      -- 
    ack_3175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 525_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_1428_inst_ack_1, ack => zeropad3D_CP_676_elements(525)); -- 
    -- CP-element group 526:  join  transition  output  bypass 
    -- CP-element group 526: predecessors 
    -- CP-element group 526: 	521 
    -- CP-element group 526: 	525 
    -- CP-element group 526: successors 
    -- CP-element group 526: 	527 
    -- CP-element group 526:  members (3) 
      -- CP-element group 526: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1431_sample_start_
      -- CP-element group 526: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1431_Sample/$entry
      -- CP-element group 526: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1431_Sample/req
      -- 
    req_3183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(526), ack => WPIPE_zeropad_output_pipe_1431_inst_req_0); -- 
    zeropad3D_cp_element_group_526: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_526"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(521) & zeropad3D_CP_676_elements(525);
      gj_zeropad3D_cp_element_group_526 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(526), clk => clk, reset => reset); --
    end block;
    -- CP-element group 527:  transition  input  output  bypass 
    -- CP-element group 527: predecessors 
    -- CP-element group 527: 	526 
    -- CP-element group 527: successors 
    -- CP-element group 527: 	528 
    -- CP-element group 527:  members (6) 
      -- CP-element group 527: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1431_sample_completed_
      -- CP-element group 527: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1431_update_start_
      -- CP-element group 527: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1431_Sample/$exit
      -- CP-element group 527: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1431_Sample/ack
      -- CP-element group 527: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1431_Update/$entry
      -- CP-element group 527: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1431_Update/req
      -- 
    ack_3184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 527_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_1431_inst_ack_0, ack => zeropad3D_CP_676_elements(527)); -- 
    req_3188_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3188_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(527), ack => WPIPE_zeropad_output_pipe_1431_inst_req_1); -- 
    -- CP-element group 528:  transition  input  bypass 
    -- CP-element group 528: predecessors 
    -- CP-element group 528: 	527 
    -- CP-element group 528: successors 
    -- CP-element group 528: 	529 
    -- CP-element group 528:  members (3) 
      -- CP-element group 528: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1431_update_completed_
      -- CP-element group 528: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1431_Update/$exit
      -- CP-element group 528: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1431_Update/ack
      -- 
    ack_3189_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 528_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_1431_inst_ack_1, ack => zeropad3D_CP_676_elements(528)); -- 
    -- CP-element group 529:  join  transition  output  bypass 
    -- CP-element group 529: predecessors 
    -- CP-element group 529: 	519 
    -- CP-element group 529: 	528 
    -- CP-element group 529: successors 
    -- CP-element group 529: 	530 
    -- CP-element group 529:  members (3) 
      -- CP-element group 529: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1434_sample_start_
      -- CP-element group 529: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1434_Sample/$entry
      -- CP-element group 529: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1434_Sample/req
      -- 
    req_3197_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3197_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(529), ack => WPIPE_zeropad_output_pipe_1434_inst_req_0); -- 
    zeropad3D_cp_element_group_529: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_529"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(519) & zeropad3D_CP_676_elements(528);
      gj_zeropad3D_cp_element_group_529 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(529), clk => clk, reset => reset); --
    end block;
    -- CP-element group 530:  transition  input  output  bypass 
    -- CP-element group 530: predecessors 
    -- CP-element group 530: 	529 
    -- CP-element group 530: successors 
    -- CP-element group 530: 	531 
    -- CP-element group 530:  members (6) 
      -- CP-element group 530: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1434_sample_completed_
      -- CP-element group 530: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1434_update_start_
      -- CP-element group 530: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1434_Sample/$exit
      -- CP-element group 530: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1434_Sample/ack
      -- CP-element group 530: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1434_Update/$entry
      -- CP-element group 530: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1434_Update/req
      -- 
    ack_3198_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 530_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_1434_inst_ack_0, ack => zeropad3D_CP_676_elements(530)); -- 
    req_3202_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3202_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(530), ack => WPIPE_zeropad_output_pipe_1434_inst_req_1); -- 
    -- CP-element group 531:  transition  input  bypass 
    -- CP-element group 531: predecessors 
    -- CP-element group 531: 	530 
    -- CP-element group 531: successors 
    -- CP-element group 531: 	532 
    -- CP-element group 531:  members (3) 
      -- CP-element group 531: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1434_update_completed_
      -- CP-element group 531: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1434_Update/$exit
      -- CP-element group 531: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1434_Update/ack
      -- 
    ack_3203_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 531_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_1434_inst_ack_1, ack => zeropad3D_CP_676_elements(531)); -- 
    -- CP-element group 532:  join  transition  output  bypass 
    -- CP-element group 532: predecessors 
    -- CP-element group 532: 	531 
    -- CP-element group 532: 	517 
    -- CP-element group 532: successors 
    -- CP-element group 532: 	533 
    -- CP-element group 532:  members (3) 
      -- CP-element group 532: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1437_sample_start_
      -- CP-element group 532: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1437_Sample/$entry
      -- CP-element group 532: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1437_Sample/req
      -- 
    req_3211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(532), ack => WPIPE_zeropad_output_pipe_1437_inst_req_0); -- 
    zeropad3D_cp_element_group_532: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_532"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(531) & zeropad3D_CP_676_elements(517);
      gj_zeropad3D_cp_element_group_532 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(532), clk => clk, reset => reset); --
    end block;
    -- CP-element group 533:  transition  input  output  bypass 
    -- CP-element group 533: predecessors 
    -- CP-element group 533: 	532 
    -- CP-element group 533: successors 
    -- CP-element group 533: 	534 
    -- CP-element group 533:  members (6) 
      -- CP-element group 533: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1437_sample_completed_
      -- CP-element group 533: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1437_update_start_
      -- CP-element group 533: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1437_Sample/$exit
      -- CP-element group 533: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1437_Sample/ack
      -- CP-element group 533: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1437_Update/$entry
      -- CP-element group 533: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1437_Update/req
      -- 
    ack_3212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 533_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_1437_inst_ack_0, ack => zeropad3D_CP_676_elements(533)); -- 
    req_3216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(533), ack => WPIPE_zeropad_output_pipe_1437_inst_req_1); -- 
    -- CP-element group 534:  transition  input  bypass 
    -- CP-element group 534: predecessors 
    -- CP-element group 534: 	533 
    -- CP-element group 534: successors 
    -- CP-element group 534: 	535 
    -- CP-element group 534:  members (3) 
      -- CP-element group 534: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1437_update_completed_
      -- CP-element group 534: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1437_Update/$exit
      -- CP-element group 534: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1437_Update/ack
      -- 
    ack_3217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 534_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_1437_inst_ack_1, ack => zeropad3D_CP_676_elements(534)); -- 
    -- CP-element group 535:  join  transition  output  bypass 
    -- CP-element group 535: predecessors 
    -- CP-element group 535: 	534 
    -- CP-element group 535: 	515 
    -- CP-element group 535: successors 
    -- CP-element group 535: 	536 
    -- CP-element group 535:  members (3) 
      -- CP-element group 535: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1440_sample_start_
      -- CP-element group 535: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1440_Sample/$entry
      -- CP-element group 535: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1440_Sample/req
      -- 
    req_3225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(535), ack => WPIPE_zeropad_output_pipe_1440_inst_req_0); -- 
    zeropad3D_cp_element_group_535: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_535"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(534) & zeropad3D_CP_676_elements(515);
      gj_zeropad3D_cp_element_group_535 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(535), clk => clk, reset => reset); --
    end block;
    -- CP-element group 536:  transition  input  output  bypass 
    -- CP-element group 536: predecessors 
    -- CP-element group 536: 	535 
    -- CP-element group 536: successors 
    -- CP-element group 536: 	537 
    -- CP-element group 536:  members (6) 
      -- CP-element group 536: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1440_sample_completed_
      -- CP-element group 536: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1440_update_start_
      -- CP-element group 536: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1440_Sample/$exit
      -- CP-element group 536: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1440_Sample/ack
      -- CP-element group 536: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1440_Update/$entry
      -- CP-element group 536: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1440_Update/req
      -- 
    ack_3226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 536_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_1440_inst_ack_0, ack => zeropad3D_CP_676_elements(536)); -- 
    req_3230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(536), ack => WPIPE_zeropad_output_pipe_1440_inst_req_1); -- 
    -- CP-element group 537:  transition  input  bypass 
    -- CP-element group 537: predecessors 
    -- CP-element group 537: 	536 
    -- CP-element group 537: successors 
    -- CP-element group 537: 	538 
    -- CP-element group 537:  members (3) 
      -- CP-element group 537: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1440_update_completed_
      -- CP-element group 537: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1440_Update/$exit
      -- CP-element group 537: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1440_Update/ack
      -- 
    ack_3231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 537_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_1440_inst_ack_1, ack => zeropad3D_CP_676_elements(537)); -- 
    -- CP-element group 538:  join  transition  output  bypass 
    -- CP-element group 538: predecessors 
    -- CP-element group 538: 	513 
    -- CP-element group 538: 	537 
    -- CP-element group 538: successors 
    -- CP-element group 538: 	539 
    -- CP-element group 538:  members (3) 
      -- CP-element group 538: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1443_sample_start_
      -- CP-element group 538: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1443_Sample/$entry
      -- CP-element group 538: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1443_Sample/req
      -- 
    req_3239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(538), ack => WPIPE_zeropad_output_pipe_1443_inst_req_0); -- 
    zeropad3D_cp_element_group_538: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_538"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(513) & zeropad3D_CP_676_elements(537);
      gj_zeropad3D_cp_element_group_538 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(538), clk => clk, reset => reset); --
    end block;
    -- CP-element group 539:  transition  input  output  bypass 
    -- CP-element group 539: predecessors 
    -- CP-element group 539: 	538 
    -- CP-element group 539: successors 
    -- CP-element group 539: 	540 
    -- CP-element group 539:  members (6) 
      -- CP-element group 539: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1443_sample_completed_
      -- CP-element group 539: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1443_update_start_
      -- CP-element group 539: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1443_Sample/$exit
      -- CP-element group 539: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1443_Sample/ack
      -- CP-element group 539: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1443_Update/$entry
      -- CP-element group 539: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1443_Update/req
      -- 
    ack_3240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 539_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_1443_inst_ack_0, ack => zeropad3D_CP_676_elements(539)); -- 
    req_3244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(539), ack => WPIPE_zeropad_output_pipe_1443_inst_req_1); -- 
    -- CP-element group 540:  transition  input  bypass 
    -- CP-element group 540: predecessors 
    -- CP-element group 540: 	539 
    -- CP-element group 540: successors 
    -- CP-element group 540: 	541 
    -- CP-element group 540:  members (3) 
      -- CP-element group 540: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1443_update_completed_
      -- CP-element group 540: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1443_Update/$exit
      -- CP-element group 540: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1443_Update/ack
      -- 
    ack_3245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 540_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_1443_inst_ack_1, ack => zeropad3D_CP_676_elements(540)); -- 
    -- CP-element group 541:  join  transition  output  bypass 
    -- CP-element group 541: predecessors 
    -- CP-element group 541: 	511 
    -- CP-element group 541: 	540 
    -- CP-element group 541: successors 
    -- CP-element group 541: 	542 
    -- CP-element group 541:  members (3) 
      -- CP-element group 541: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1446_sample_start_
      -- CP-element group 541: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1446_Sample/$entry
      -- CP-element group 541: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1446_Sample/req
      -- 
    req_3253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(541), ack => WPIPE_zeropad_output_pipe_1446_inst_req_0); -- 
    zeropad3D_cp_element_group_541: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_541"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(511) & zeropad3D_CP_676_elements(540);
      gj_zeropad3D_cp_element_group_541 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(541), clk => clk, reset => reset); --
    end block;
    -- CP-element group 542:  transition  input  output  bypass 
    -- CP-element group 542: predecessors 
    -- CP-element group 542: 	541 
    -- CP-element group 542: successors 
    -- CP-element group 542: 	543 
    -- CP-element group 542:  members (6) 
      -- CP-element group 542: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1446_sample_completed_
      -- CP-element group 542: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1446_update_start_
      -- CP-element group 542: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1446_Sample/$exit
      -- CP-element group 542: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1446_Sample/ack
      -- CP-element group 542: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1446_Update/$entry
      -- CP-element group 542: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1446_Update/req
      -- 
    ack_3254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 542_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_1446_inst_ack_0, ack => zeropad3D_CP_676_elements(542)); -- 
    req_3258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(542), ack => WPIPE_zeropad_output_pipe_1446_inst_req_1); -- 
    -- CP-element group 543:  transition  input  bypass 
    -- CP-element group 543: predecessors 
    -- CP-element group 543: 	542 
    -- CP-element group 543: successors 
    -- CP-element group 543: 	544 
    -- CP-element group 543:  members (3) 
      -- CP-element group 543: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1446_update_completed_
      -- CP-element group 543: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1446_Update/$exit
      -- CP-element group 543: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1446_Update/ack
      -- 
    ack_3259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 543_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_1446_inst_ack_1, ack => zeropad3D_CP_676_elements(543)); -- 
    -- CP-element group 544:  join  transition  output  bypass 
    -- CP-element group 544: predecessors 
    -- CP-element group 544: 	543 
    -- CP-element group 544: 	509 
    -- CP-element group 544: successors 
    -- CP-element group 544: 	545 
    -- CP-element group 544:  members (3) 
      -- CP-element group 544: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1449_sample_start_
      -- CP-element group 544: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1449_Sample/$entry
      -- CP-element group 544: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1449_Sample/req
      -- 
    req_3267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(544), ack => WPIPE_zeropad_output_pipe_1449_inst_req_0); -- 
    zeropad3D_cp_element_group_544: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_544"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(543) & zeropad3D_CP_676_elements(509);
      gj_zeropad3D_cp_element_group_544 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(544), clk => clk, reset => reset); --
    end block;
    -- CP-element group 545:  transition  input  output  bypass 
    -- CP-element group 545: predecessors 
    -- CP-element group 545: 	544 
    -- CP-element group 545: successors 
    -- CP-element group 545: 	546 
    -- CP-element group 545:  members (6) 
      -- CP-element group 545: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1449_sample_completed_
      -- CP-element group 545: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1449_update_start_
      -- CP-element group 545: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1449_Sample/$exit
      -- CP-element group 545: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1449_Sample/ack
      -- CP-element group 545: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1449_Update/$entry
      -- CP-element group 545: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1449_Update/req
      -- 
    ack_3268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 545_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_1449_inst_ack_0, ack => zeropad3D_CP_676_elements(545)); -- 
    req_3272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(545), ack => WPIPE_zeropad_output_pipe_1449_inst_req_1); -- 
    -- CP-element group 546:  fork  transition  place  input  output  bypass 
    -- CP-element group 546: predecessors 
    -- CP-element group 546: 	545 
    -- CP-element group 546: successors 
    -- CP-element group 546: 	547 
    -- CP-element group 546: 	548 
    -- CP-element group 546: 	549 
    -- CP-element group 546: 	550 
    -- CP-element group 546: 	553 
    -- CP-element group 546:  members (22) 
      -- CP-element group 546: 	 branch_block_stmt_222/assign_stmt_1456_to_call_stmt_1472__entry__
      -- CP-element group 546: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451__exit__
      -- CP-element group 546: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/$exit
      -- CP-element group 546: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1449_update_completed_
      -- CP-element group 546: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1449_Update/$exit
      -- CP-element group 546: 	 branch_block_stmt_222/call_stmt_1343_to_assign_stmt_1451/WPIPE_zeropad_output_pipe_1449_Update/ack
      -- CP-element group 546: 	 branch_block_stmt_222/assign_stmt_1456_to_call_stmt_1472/$entry
      -- CP-element group 546: 	 branch_block_stmt_222/assign_stmt_1456_to_call_stmt_1472/type_cast_1455_sample_start_
      -- CP-element group 546: 	 branch_block_stmt_222/assign_stmt_1456_to_call_stmt_1472/type_cast_1455_update_start_
      -- CP-element group 546: 	 branch_block_stmt_222/assign_stmt_1456_to_call_stmt_1472/type_cast_1455_Sample/$entry
      -- CP-element group 546: 	 branch_block_stmt_222/assign_stmt_1456_to_call_stmt_1472/type_cast_1455_Sample/rr
      -- CP-element group 546: 	 branch_block_stmt_222/assign_stmt_1456_to_call_stmt_1472/type_cast_1455_Update/$entry
      -- CP-element group 546: 	 branch_block_stmt_222/assign_stmt_1456_to_call_stmt_1472/type_cast_1455_Update/cr
      -- CP-element group 546: 	 branch_block_stmt_222/assign_stmt_1456_to_call_stmt_1472/type_cast_1459_sample_start_
      -- CP-element group 546: 	 branch_block_stmt_222/assign_stmt_1456_to_call_stmt_1472/type_cast_1459_update_start_
      -- CP-element group 546: 	 branch_block_stmt_222/assign_stmt_1456_to_call_stmt_1472/type_cast_1459_Sample/$entry
      -- CP-element group 546: 	 branch_block_stmt_222/assign_stmt_1456_to_call_stmt_1472/type_cast_1459_Sample/rr
      -- CP-element group 546: 	 branch_block_stmt_222/assign_stmt_1456_to_call_stmt_1472/type_cast_1459_Update/$entry
      -- CP-element group 546: 	 branch_block_stmt_222/assign_stmt_1456_to_call_stmt_1472/type_cast_1459_Update/cr
      -- CP-element group 546: 	 branch_block_stmt_222/assign_stmt_1456_to_call_stmt_1472/call_stmt_1472_update_start_
      -- CP-element group 546: 	 branch_block_stmt_222/assign_stmt_1456_to_call_stmt_1472/call_stmt_1472_Update/$entry
      -- CP-element group 546: 	 branch_block_stmt_222/assign_stmt_1456_to_call_stmt_1472/call_stmt_1472_Update/ccr
      -- 
    ack_3273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 546_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_1449_inst_ack_1, ack => zeropad3D_CP_676_elements(546)); -- 
    rr_3284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(546), ack => type_cast_1455_inst_req_0); -- 
    cr_3289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(546), ack => type_cast_1455_inst_req_1); -- 
    rr_3298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(546), ack => type_cast_1459_inst_req_0); -- 
    cr_3303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(546), ack => type_cast_1459_inst_req_1); -- 
    ccr_3317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(546), ack => call_stmt_1472_call_req_1); -- 
    -- CP-element group 547:  transition  input  bypass 
    -- CP-element group 547: predecessors 
    -- CP-element group 547: 	546 
    -- CP-element group 547: successors 
    -- CP-element group 547:  members (3) 
      -- CP-element group 547: 	 branch_block_stmt_222/assign_stmt_1456_to_call_stmt_1472/type_cast_1455_sample_completed_
      -- CP-element group 547: 	 branch_block_stmt_222/assign_stmt_1456_to_call_stmt_1472/type_cast_1455_Sample/$exit
      -- CP-element group 547: 	 branch_block_stmt_222/assign_stmt_1456_to_call_stmt_1472/type_cast_1455_Sample/ra
      -- 
    ra_3285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 547_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1455_inst_ack_0, ack => zeropad3D_CP_676_elements(547)); -- 
    -- CP-element group 548:  transition  input  bypass 
    -- CP-element group 548: predecessors 
    -- CP-element group 548: 	546 
    -- CP-element group 548: successors 
    -- CP-element group 548: 	551 
    -- CP-element group 548:  members (3) 
      -- CP-element group 548: 	 branch_block_stmt_222/assign_stmt_1456_to_call_stmt_1472/type_cast_1455_update_completed_
      -- CP-element group 548: 	 branch_block_stmt_222/assign_stmt_1456_to_call_stmt_1472/type_cast_1455_Update/$exit
      -- CP-element group 548: 	 branch_block_stmt_222/assign_stmt_1456_to_call_stmt_1472/type_cast_1455_Update/ca
      -- 
    ca_3290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 548_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1455_inst_ack_1, ack => zeropad3D_CP_676_elements(548)); -- 
    -- CP-element group 549:  transition  input  bypass 
    -- CP-element group 549: predecessors 
    -- CP-element group 549: 	546 
    -- CP-element group 549: successors 
    -- CP-element group 549:  members (3) 
      -- CP-element group 549: 	 branch_block_stmt_222/assign_stmt_1456_to_call_stmt_1472/type_cast_1459_sample_completed_
      -- CP-element group 549: 	 branch_block_stmt_222/assign_stmt_1456_to_call_stmt_1472/type_cast_1459_Sample/$exit
      -- CP-element group 549: 	 branch_block_stmt_222/assign_stmt_1456_to_call_stmt_1472/type_cast_1459_Sample/ra
      -- 
    ra_3299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 549_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1459_inst_ack_0, ack => zeropad3D_CP_676_elements(549)); -- 
    -- CP-element group 550:  transition  input  bypass 
    -- CP-element group 550: predecessors 
    -- CP-element group 550: 	546 
    -- CP-element group 550: successors 
    -- CP-element group 550: 	551 
    -- CP-element group 550:  members (3) 
      -- CP-element group 550: 	 branch_block_stmt_222/assign_stmt_1456_to_call_stmt_1472/type_cast_1459_update_completed_
      -- CP-element group 550: 	 branch_block_stmt_222/assign_stmt_1456_to_call_stmt_1472/type_cast_1459_Update/$exit
      -- CP-element group 550: 	 branch_block_stmt_222/assign_stmt_1456_to_call_stmt_1472/type_cast_1459_Update/ca
      -- 
    ca_3304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 550_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1459_inst_ack_1, ack => zeropad3D_CP_676_elements(550)); -- 
    -- CP-element group 551:  join  transition  output  bypass 
    -- CP-element group 551: predecessors 
    -- CP-element group 551: 	548 
    -- CP-element group 551: 	550 
    -- CP-element group 551: successors 
    -- CP-element group 551: 	552 
    -- CP-element group 551:  members (3) 
      -- CP-element group 551: 	 branch_block_stmt_222/assign_stmt_1456_to_call_stmt_1472/call_stmt_1472_sample_start_
      -- CP-element group 551: 	 branch_block_stmt_222/assign_stmt_1456_to_call_stmt_1472/call_stmt_1472_Sample/$entry
      -- CP-element group 551: 	 branch_block_stmt_222/assign_stmt_1456_to_call_stmt_1472/call_stmt_1472_Sample/crr
      -- 
    crr_3312_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3312_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(551), ack => call_stmt_1472_call_req_0); -- 
    zeropad3D_cp_element_group_551: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_551"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(548) & zeropad3D_CP_676_elements(550);
      gj_zeropad3D_cp_element_group_551 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(551), clk => clk, reset => reset); --
    end block;
    -- CP-element group 552:  transition  input  bypass 
    -- CP-element group 552: predecessors 
    -- CP-element group 552: 	551 
    -- CP-element group 552: successors 
    -- CP-element group 552:  members (3) 
      -- CP-element group 552: 	 branch_block_stmt_222/assign_stmt_1456_to_call_stmt_1472/call_stmt_1472_sample_completed_
      -- CP-element group 552: 	 branch_block_stmt_222/assign_stmt_1456_to_call_stmt_1472/call_stmt_1472_Sample/$exit
      -- CP-element group 552: 	 branch_block_stmt_222/assign_stmt_1456_to_call_stmt_1472/call_stmt_1472_Sample/cra
      -- 
    cra_3313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 552_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1472_call_ack_0, ack => zeropad3D_CP_676_elements(552)); -- 
    -- CP-element group 553:  transition  place  input  bypass 
    -- CP-element group 553: predecessors 
    -- CP-element group 553: 	546 
    -- CP-element group 553: successors 
    -- CP-element group 553:  members (16) 
      -- CP-element group 553: 	 branch_block_stmt_222/merge_stmt_1474__exit__
      -- CP-element group 553: 	 branch_block_stmt_222/return__
      -- CP-element group 553: 	 branch_block_stmt_222/assign_stmt_1456_to_call_stmt_1472__exit__
      -- CP-element group 553: 	 branch_block_stmt_222/branch_block_stmt_222__exit__
      -- CP-element group 553: 	 branch_block_stmt_222/$exit
      -- CP-element group 553: 	 $exit
      -- CP-element group 553: 	 branch_block_stmt_222/assign_stmt_1456_to_call_stmt_1472/$exit
      -- CP-element group 553: 	 branch_block_stmt_222/assign_stmt_1456_to_call_stmt_1472/call_stmt_1472_update_completed_
      -- CP-element group 553: 	 branch_block_stmt_222/assign_stmt_1456_to_call_stmt_1472/call_stmt_1472_Update/$exit
      -- CP-element group 553: 	 branch_block_stmt_222/assign_stmt_1456_to_call_stmt_1472/call_stmt_1472_Update/cca
      -- CP-element group 553: 	 branch_block_stmt_222/return___PhiReq/$entry
      -- CP-element group 553: 	 branch_block_stmt_222/return___PhiReq/$exit
      -- CP-element group 553: 	 branch_block_stmt_222/merge_stmt_1474_PhiReqMerge
      -- CP-element group 553: 	 branch_block_stmt_222/merge_stmt_1474_PhiAck/$entry
      -- CP-element group 553: 	 branch_block_stmt_222/merge_stmt_1474_PhiAck/$exit
      -- CP-element group 553: 	 branch_block_stmt_222/merge_stmt_1474_PhiAck/dummy
      -- 
    cca_3318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 553_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1472_call_ack_1, ack => zeropad3D_CP_676_elements(553)); -- 
    -- CP-element group 554:  transition  output  delay-element  bypass 
    -- CP-element group 554: predecessors 
    -- CP-element group 554: 	70 
    -- CP-element group 554: successors 
    -- CP-element group 554: 	558 
    -- CP-element group 554:  members (5) 
      -- CP-element group 554: 	 branch_block_stmt_222/bbx_xnph_forx_xbody_PhiReq/$exit
      -- CP-element group 554: 	 branch_block_stmt_222/bbx_xnph_forx_xbody_PhiReq/phi_stmt_461/$exit
      -- CP-element group 554: 	 branch_block_stmt_222/bbx_xnph_forx_xbody_PhiReq/phi_stmt_461/phi_stmt_461_sources/$exit
      -- CP-element group 554: 	 branch_block_stmt_222/bbx_xnph_forx_xbody_PhiReq/phi_stmt_461/phi_stmt_461_sources/type_cast_465_konst_delay_trans
      -- CP-element group 554: 	 branch_block_stmt_222/bbx_xnph_forx_xbody_PhiReq/phi_stmt_461/phi_stmt_461_req
      -- 
    phi_stmt_461_req_3341_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_461_req_3341_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(554), ack => phi_stmt_461_req_0); -- 
    -- Element group zeropad3D_CP_676_elements(554) is a control-delay.
    cp_element_554_delay: control_delay_element  generic map(name => " 554_delay", delay_value => 1)  port map(req => zeropad3D_CP_676_elements(70), ack => zeropad3D_CP_676_elements(554), clk => clk, reset =>reset);
    -- CP-element group 555:  transition  input  bypass 
    -- CP-element group 555: predecessors 
    -- CP-element group 555: 	113 
    -- CP-element group 555: successors 
    -- CP-element group 555: 	557 
    -- CP-element group 555:  members (2) 
      -- CP-element group 555: 	 branch_block_stmt_222/forx_xbody_forx_xbody_PhiReq/phi_stmt_461/phi_stmt_461_sources/type_cast_467/SplitProtocol/Sample/$exit
      -- CP-element group 555: 	 branch_block_stmt_222/forx_xbody_forx_xbody_PhiReq/phi_stmt_461/phi_stmt_461_sources/type_cast_467/SplitProtocol/Sample/ra
      -- 
    ra_3361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 555_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_467_inst_ack_0, ack => zeropad3D_CP_676_elements(555)); -- 
    -- CP-element group 556:  transition  input  bypass 
    -- CP-element group 556: predecessors 
    -- CP-element group 556: 	113 
    -- CP-element group 556: successors 
    -- CP-element group 556: 	557 
    -- CP-element group 556:  members (2) 
      -- CP-element group 556: 	 branch_block_stmt_222/forx_xbody_forx_xbody_PhiReq/phi_stmt_461/phi_stmt_461_sources/type_cast_467/SplitProtocol/Update/$exit
      -- CP-element group 556: 	 branch_block_stmt_222/forx_xbody_forx_xbody_PhiReq/phi_stmt_461/phi_stmt_461_sources/type_cast_467/SplitProtocol/Update/ca
      -- 
    ca_3366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 556_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_467_inst_ack_1, ack => zeropad3D_CP_676_elements(556)); -- 
    -- CP-element group 557:  join  transition  output  bypass 
    -- CP-element group 557: predecessors 
    -- CP-element group 557: 	555 
    -- CP-element group 557: 	556 
    -- CP-element group 557: successors 
    -- CP-element group 557: 	558 
    -- CP-element group 557:  members (6) 
      -- CP-element group 557: 	 branch_block_stmt_222/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 557: 	 branch_block_stmt_222/forx_xbody_forx_xbody_PhiReq/phi_stmt_461/$exit
      -- CP-element group 557: 	 branch_block_stmt_222/forx_xbody_forx_xbody_PhiReq/phi_stmt_461/phi_stmt_461_sources/$exit
      -- CP-element group 557: 	 branch_block_stmt_222/forx_xbody_forx_xbody_PhiReq/phi_stmt_461/phi_stmt_461_sources/type_cast_467/$exit
      -- CP-element group 557: 	 branch_block_stmt_222/forx_xbody_forx_xbody_PhiReq/phi_stmt_461/phi_stmt_461_sources/type_cast_467/SplitProtocol/$exit
      -- CP-element group 557: 	 branch_block_stmt_222/forx_xbody_forx_xbody_PhiReq/phi_stmt_461/phi_stmt_461_req
      -- 
    phi_stmt_461_req_3367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_461_req_3367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(557), ack => phi_stmt_461_req_1); -- 
    zeropad3D_cp_element_group_557: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_557"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(555) & zeropad3D_CP_676_elements(556);
      gj_zeropad3D_cp_element_group_557 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(557), clk => clk, reset => reset); --
    end block;
    -- CP-element group 558:  merge  transition  place  bypass 
    -- CP-element group 558: predecessors 
    -- CP-element group 558: 	557 
    -- CP-element group 558: 	554 
    -- CP-element group 558: successors 
    -- CP-element group 558: 	559 
    -- CP-element group 558:  members (2) 
      -- CP-element group 558: 	 branch_block_stmt_222/merge_stmt_460_PhiReqMerge
      -- CP-element group 558: 	 branch_block_stmt_222/merge_stmt_460_PhiAck/$entry
      -- 
    zeropad3D_CP_676_elements(558) <= OrReduce(zeropad3D_CP_676_elements(557) & zeropad3D_CP_676_elements(554));
    -- CP-element group 559:  fork  transition  place  input  output  bypass 
    -- CP-element group 559: predecessors 
    -- CP-element group 559: 	558 
    -- CP-element group 559: successors 
    -- CP-element group 559: 	79 
    -- CP-element group 559: 	76 
    -- CP-element group 559: 	91 
    -- CP-element group 559: 	95 
    -- CP-element group 559: 	87 
    -- CP-element group 559: 	83 
    -- CP-element group 559: 	72 
    -- CP-element group 559: 	73 
    -- CP-element group 559: 	75 
    -- CP-element group 559: 	99 
    -- CP-element group 559: 	103 
    -- CP-element group 559: 	107 
    -- CP-element group 559: 	110 
    -- CP-element group 559:  members (56) 
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/ptr_deref_610_Update/word_access_complete/$entry
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/ptr_deref_610_Update/word_access_complete/word_0/cr
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623__entry__
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/ptr_deref_610_Update/word_access_complete/word_0/$entry
      -- CP-element group 559: 	 branch_block_stmt_222/merge_stmt_460__exit__
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/ptr_deref_610_Update/$entry
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/$entry
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/addr_of_474_update_start_
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/array_obj_ref_473_index_resized_1
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/array_obj_ref_473_index_scaled_1
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/array_obj_ref_473_index_computed_1
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/array_obj_ref_473_index_resize_1/$entry
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/array_obj_ref_473_index_resize_1/$exit
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/array_obj_ref_473_index_resize_1/index_resize_req
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/array_obj_ref_473_index_resize_1/index_resize_ack
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/array_obj_ref_473_index_scale_1/$entry
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/array_obj_ref_473_index_scale_1/$exit
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/array_obj_ref_473_index_scale_1/scale_rename_req
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/array_obj_ref_473_index_scale_1/scale_rename_ack
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/array_obj_ref_473_final_index_sum_regn_update_start
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/array_obj_ref_473_final_index_sum_regn_Sample/$entry
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/array_obj_ref_473_final_index_sum_regn_Sample/req
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/array_obj_ref_473_final_index_sum_regn_Update/$entry
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/array_obj_ref_473_final_index_sum_regn_Update/req
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/addr_of_474_complete/$entry
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/addr_of_474_complete/req
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_477_sample_start_
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_477_Sample/$entry
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/RPIPE_zeropad_input_pipe_477_Sample/rr
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_481_update_start_
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_481_Update/$entry
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_481_Update/cr
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_494_update_start_
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_494_Update/$entry
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_494_Update/cr
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_512_update_start_
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_512_Update/$entry
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_512_Update/cr
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_530_update_start_
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_530_Update/$entry
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_530_Update/cr
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_548_update_start_
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_548_Update/$entry
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_548_Update/cr
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_566_update_start_
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_566_Update/$entry
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_566_Update/cr
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_584_update_start_
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_584_Update/$entry
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_584_Update/cr
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_602_update_start_
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_602_Update/$entry
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/type_cast_602_Update/cr
      -- CP-element group 559: 	 branch_block_stmt_222/assign_stmt_475_to_assign_stmt_623/ptr_deref_610_update_start_
      -- CP-element group 559: 	 branch_block_stmt_222/merge_stmt_460_PhiAck/$exit
      -- CP-element group 559: 	 branch_block_stmt_222/merge_stmt_460_PhiAck/phi_stmt_461_ack
      -- 
    phi_stmt_461_ack_3372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 559_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_461_ack_0, ack => zeropad3D_CP_676_elements(559)); -- 
    cr_1514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(559), ack => ptr_deref_610_store_0_req_1); -- 
    req_1220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(559), ack => array_obj_ref_473_index_offset_req_0); -- 
    req_1225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(559), ack => array_obj_ref_473_index_offset_req_1); -- 
    req_1240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(559), ack => addr_of_474_final_reg_req_1); -- 
    rr_1249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(559), ack => RPIPE_zeropad_input_pipe_477_inst_req_0); -- 
    cr_1268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(559), ack => type_cast_481_inst_req_1); -- 
    cr_1296_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1296_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(559), ack => type_cast_494_inst_req_1); -- 
    cr_1324_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1324_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(559), ack => type_cast_512_inst_req_1); -- 
    cr_1352_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1352_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(559), ack => type_cast_530_inst_req_1); -- 
    cr_1380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(559), ack => type_cast_548_inst_req_1); -- 
    cr_1408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(559), ack => type_cast_566_inst_req_1); -- 
    cr_1436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(559), ack => type_cast_584_inst_req_1); -- 
    cr_1464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(559), ack => type_cast_602_inst_req_1); -- 
    -- CP-element group 560:  merge  fork  transition  place  output  bypass 
    -- CP-element group 560: predecessors 
    -- CP-element group 560: 	71 
    -- CP-element group 560: 	112 
    -- CP-element group 560: successors 
    -- CP-element group 560: 	114 
    -- CP-element group 560: 	115 
    -- CP-element group 560: 	116 
    -- CP-element group 560: 	117 
    -- CP-element group 560: 	118 
    -- CP-element group 560: 	119 
    -- CP-element group 560: 	120 
    -- CP-element group 560: 	121 
    -- CP-element group 560: 	122 
    -- CP-element group 560: 	123 
    -- CP-element group 560: 	124 
    -- CP-element group 560: 	125 
    -- CP-element group 560:  members (43) 
      -- CP-element group 560: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_649_Sample/$entry
      -- CP-element group 560: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_653_Update/cr
      -- CP-element group 560: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688__entry__
      -- CP-element group 560: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_649_update_start_
      -- CP-element group 560: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_649_Sample/rr
      -- CP-element group 560: 	 branch_block_stmt_222/merge_stmt_632__exit__
      -- CP-element group 560: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_649_Update/$entry
      -- CP-element group 560: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_645_Update/cr
      -- CP-element group 560: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_653_sample_start_
      -- CP-element group 560: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_649_Update/cr
      -- CP-element group 560: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_653_update_start_
      -- CP-element group 560: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_649_sample_start_
      -- CP-element group 560: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_668_update_start_
      -- CP-element group 560: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_653_Sample/$entry
      -- CP-element group 560: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_645_Sample/rr
      -- CP-element group 560: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_645_Update/$entry
      -- CP-element group 560: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_645_Sample/$entry
      -- CP-element group 560: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_645_update_start_
      -- CP-element group 560: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_653_Update/$entry
      -- CP-element group 560: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_653_Sample/rr
      -- CP-element group 560: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_645_sample_start_
      -- CP-element group 560: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/call_stmt_635_Update/ccr
      -- CP-element group 560: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_668_sample_start_
      -- CP-element group 560: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/call_stmt_635_Update/$entry
      -- CP-element group 560: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/call_stmt_635_Sample/crr
      -- CP-element group 560: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/call_stmt_635_Sample/$entry
      -- CP-element group 560: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/call_stmt_635_update_start_
      -- CP-element group 560: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/call_stmt_635_sample_start_
      -- CP-element group 560: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/$entry
      -- CP-element group 560: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_677_Update/cr
      -- CP-element group 560: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_677_Update/$entry
      -- CP-element group 560: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_677_Sample/rr
      -- CP-element group 560: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_677_Sample/$entry
      -- CP-element group 560: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_677_update_start_
      -- CP-element group 560: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_677_sample_start_
      -- CP-element group 560: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_668_Update/cr
      -- CP-element group 560: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_668_Update/$entry
      -- CP-element group 560: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_668_Sample/rr
      -- CP-element group 560: 	 branch_block_stmt_222/call_stmt_635_to_assign_stmt_688/type_cast_668_Sample/$entry
      -- CP-element group 560: 	 branch_block_stmt_222/merge_stmt_632_PhiReqMerge
      -- CP-element group 560: 	 branch_block_stmt_222/merge_stmt_632_PhiAck/$entry
      -- CP-element group 560: 	 branch_block_stmt_222/merge_stmt_632_PhiAck/$exit
      -- CP-element group 560: 	 branch_block_stmt_222/merge_stmt_632_PhiAck/dummy
      -- 
    cr_1592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(560), ack => type_cast_653_inst_req_1); -- 
    rr_1573_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1573_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(560), ack => type_cast_649_inst_req_0); -- 
    cr_1564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(560), ack => type_cast_645_inst_req_1); -- 
    cr_1578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(560), ack => type_cast_649_inst_req_1); -- 
    rr_1559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(560), ack => type_cast_645_inst_req_0); -- 
    rr_1587_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1587_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(560), ack => type_cast_653_inst_req_0); -- 
    ccr_1550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(560), ack => call_stmt_635_call_req_1); -- 
    crr_1545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(560), ack => call_stmt_635_call_req_0); -- 
    cr_1620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(560), ack => type_cast_677_inst_req_1); -- 
    rr_1615_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1615_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(560), ack => type_cast_677_inst_req_0); -- 
    cr_1606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(560), ack => type_cast_668_inst_req_1); -- 
    rr_1601_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1601_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(560), ack => type_cast_668_inst_req_0); -- 
    zeropad3D_CP_676_elements(560) <= OrReduce(zeropad3D_CP_676_elements(71) & zeropad3D_CP_676_elements(112));
    zeropad3D_do_while_stmt_707_terminator_2983: loop_terminator -- 
      generic map (name => " zeropad3D_do_while_stmt_707_terminator_2983", max_iterations_in_flight =>15) 
      port map(loop_body_exit => zeropad3D_CP_676_elements(131),loop_continue => zeropad3D_CP_676_elements(498),loop_terminate => zeropad3D_CP_676_elements(497),loop_back => zeropad3D_CP_676_elements(129),loop_exit => zeropad3D_CP_676_elements(128),clk => clk, reset => reset); -- 
    phi_stmt_709_phi_seq_1685_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= zeropad3D_CP_676_elements(144);
      zeropad3D_CP_676_elements(149)<= src_sample_reqs(0);
      src_sample_acks(0)  <= zeropad3D_CP_676_elements(153);
      zeropad3D_CP_676_elements(150)<= src_update_reqs(0);
      src_update_acks(0)  <= zeropad3D_CP_676_elements(154);
      zeropad3D_CP_676_elements(145) <= phi_mux_reqs(0);
      triggers(1)  <= zeropad3D_CP_676_elements(146);
      zeropad3D_CP_676_elements(155)<= src_sample_reqs(1);
      src_sample_acks(1)  <= zeropad3D_CP_676_elements(155);
      zeropad3D_CP_676_elements(156)<= src_update_reqs(1);
      src_update_acks(1)  <= zeropad3D_CP_676_elements(157);
      zeropad3D_CP_676_elements(147) <= phi_mux_reqs(1);
      phi_stmt_709_phi_seq_1685 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_709_phi_seq_1685") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => zeropad3D_CP_676_elements(136), 
          phi_sample_ack => zeropad3D_CP_676_elements(142), 
          phi_update_req => zeropad3D_CP_676_elements(138), 
          phi_update_ack => zeropad3D_CP_676_elements(143), 
          phi_mux_ack => zeropad3D_CP_676_elements(148), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_714_phi_seq_1729_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= zeropad3D_CP_676_elements(165);
      zeropad3D_CP_676_elements(170)<= src_sample_reqs(0);
      src_sample_acks(0)  <= zeropad3D_CP_676_elements(174);
      zeropad3D_CP_676_elements(171)<= src_update_reqs(0);
      src_update_acks(0)  <= zeropad3D_CP_676_elements(175);
      zeropad3D_CP_676_elements(166) <= phi_mux_reqs(0);
      triggers(1)  <= zeropad3D_CP_676_elements(167);
      zeropad3D_CP_676_elements(176)<= src_sample_reqs(1);
      src_sample_acks(1)  <= zeropad3D_CP_676_elements(176);
      zeropad3D_CP_676_elements(177)<= src_update_reqs(1);
      src_update_acks(1)  <= zeropad3D_CP_676_elements(178);
      zeropad3D_CP_676_elements(168) <= phi_mux_reqs(1);
      phi_stmt_714_phi_seq_1729 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_714_phi_seq_1729") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => zeropad3D_CP_676_elements(161), 
          phi_sample_ack => zeropad3D_CP_676_elements(162), 
          phi_update_req => zeropad3D_CP_676_elements(163), 
          phi_update_ack => zeropad3D_CP_676_elements(164), 
          phi_mux_ack => zeropad3D_CP_676_elements(169), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_719_phi_seq_1773_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= zeropad3D_CP_676_elements(186);
      zeropad3D_CP_676_elements(191)<= src_sample_reqs(0);
      src_sample_acks(0)  <= zeropad3D_CP_676_elements(195);
      zeropad3D_CP_676_elements(192)<= src_update_reqs(0);
      src_update_acks(0)  <= zeropad3D_CP_676_elements(196);
      zeropad3D_CP_676_elements(187) <= phi_mux_reqs(0);
      triggers(1)  <= zeropad3D_CP_676_elements(188);
      zeropad3D_CP_676_elements(197)<= src_sample_reqs(1);
      src_sample_acks(1)  <= zeropad3D_CP_676_elements(197);
      zeropad3D_CP_676_elements(198)<= src_update_reqs(1);
      src_update_acks(1)  <= zeropad3D_CP_676_elements(199);
      zeropad3D_CP_676_elements(189) <= phi_mux_reqs(1);
      phi_stmt_719_phi_seq_1773 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_719_phi_seq_1773") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => zeropad3D_CP_676_elements(182), 
          phi_sample_ack => zeropad3D_CP_676_elements(183), 
          phi_update_req => zeropad3D_CP_676_elements(184), 
          phi_update_ack => zeropad3D_CP_676_elements(185), 
          phi_mux_ack => zeropad3D_CP_676_elements(190), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1637_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= zeropad3D_CP_676_elements(132);
        preds(1)  <= zeropad3D_CP_676_elements(133);
        entry_tmerge_1637 : transition_merge -- 
          generic map(name => " entry_tmerge_1637")
          port map (preds => preds, symbol_out => zeropad3D_CP_676_elements(134));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_1196_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1243_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1289_wire : std_logic_vector(31 downto 0);
    signal ASHR_i64_i64_424_wire : std_logic_vector(63 downto 0);
    signal MUX_893_wire : std_logic_vector(15 downto 0);
    signal MUX_894_wire : std_logic_vector(15 downto 0);
    signal MUX_921_wire : std_logic_vector(15 downto 0);
    signal MUX_922_wire : std_logic_vector(15 downto 0);
    signal MUX_949_wire : std_logic_vector(15 downto 0);
    signal MUX_950_wire : std_logic_vector(15 downto 0);
    signal MUX_971_wire : std_logic_vector(15 downto 0);
    signal MUX_972_wire : std_logic_vector(15 downto 0);
    signal NOT_u1_u1_1096_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1166_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_854_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_870_wire : std_logic_vector(0 downto 0);
    signal R_idxprom290_1211_resized : std_logic_vector(13 downto 0);
    signal R_idxprom290_1211_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom296_1258_resized : std_logic_vector(13 downto 0);
    signal R_idxprom296_1258_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom302_1304_resized : std_logic_vector(13 downto 0);
    signal R_idxprom302_1304_scaled : std_logic_vector(13 downto 0);
    signal R_indvar_472_resized : std_logic_vector(13 downto 0);
    signal R_indvar_472_scaled : std_logic_vector(13 downto 0);
    signal add104_536 : std_logic_vector(63 downto 0);
    signal add110_554 : std_logic_vector(63 downto 0);
    signal add116_572 : std_logic_vector(63 downto 0);
    signal add122_590 : std_logic_vector(63 downto 0);
    signal add128_608 : std_logic_vector(63 downto 0);
    signal add184_758 : std_logic_vector(15 downto 0);
    signal add195_665 : std_logic_vector(31 downto 0);
    signal add209_674 : std_logic_vector(31 downto 0);
    signal add230_1056_delayed_2_0_1179 : std_logic_vector(15 downto 0);
    signal add230_1128_delayed_2_0_1272 : std_logic_vector(15 downto 0);
    signal add230_998 : std_logic_vector(15 downto 0);
    signal add23_260 : std_logic_vector(15 downto 0);
    signal add252_1034 : std_logic_vector(15 downto 0);
    signal add252_1094_delayed_2_0_1226 : std_logic_vector(15 downto 0);
    signal add266_683 : std_logic_vector(31 downto 0);
    signal add283_688 : std_logic_vector(31 downto 0);
    signal add32_285 : std_logic_vector(15 downto 0);
    signal add41_310 : std_logic_vector(15 downto 0);
    signal add51_338 : std_logic_vector(31 downto 0);
    signal add60_363 : std_logic_vector(15 downto 0);
    signal add69_388 : std_logic_vector(15 downto 0);
    signal add92_500 : std_logic_vector(63 downto 0);
    signal add98_518 : std_logic_vector(63 downto 0);
    signal array_obj_ref_1212_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1212_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1212_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1212_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1212_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1212_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1259_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1259_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1259_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1259_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1259_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1259_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1305_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1305_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1305_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1305_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1305_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1305_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_473_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_473_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_473_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_473_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_473_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_473_root_address : std_logic_vector(13 downto 0);
    signal arrayidx291_1214 : std_logic_vector(31 downto 0);
    signal arrayidx297_1261 : std_logic_vector(31 downto 0);
    signal arrayidx303_1156_delayed_5_0_1313 : std_logic_vector(31 downto 0);
    signal arrayidx303_1307 : std_logic_vector(31 downto 0);
    signal arrayidx_475 : std_logic_vector(31 downto 0);
    signal call101_527 : std_logic_vector(7 downto 0);
    signal call107_545 : std_logic_vector(7 downto 0);
    signal call113_563 : std_logic_vector(7 downto 0);
    signal call119_581 : std_logic_vector(7 downto 0);
    signal call11_234 : std_logic_vector(7 downto 0);
    signal call125_599 : std_logic_vector(7 downto 0);
    signal call133_635 : std_logic_vector(63 downto 0);
    signal call16_237 : std_logic_vector(7 downto 0);
    signal call21_251 : std_logic_vector(7 downto 0);
    signal call25_263 : std_logic_vector(7 downto 0);
    signal call2_228 : std_logic_vector(7 downto 0);
    signal call309_1343 : std_logic_vector(63 downto 0);
    signal call30_276 : std_logic_vector(7 downto 0);
    signal call34_288 : std_logic_vector(7 downto 0);
    signal call39_301 : std_logic_vector(7 downto 0);
    signal call43_313 : std_logic_vector(7 downto 0);
    signal call44_316 : std_logic_vector(7 downto 0);
    signal call49_329 : std_logic_vector(7 downto 0);
    signal call53_341 : std_logic_vector(7 downto 0);
    signal call58_354 : std_logic_vector(7 downto 0);
    signal call62_366 : std_logic_vector(7 downto 0);
    signal call67_379 : std_logic_vector(7 downto 0);
    signal call6_231 : std_logic_vector(7 downto 0);
    signal call85_478 : std_logic_vector(7 downto 0);
    signal call89_491 : std_logic_vector(7 downto 0);
    signal call95_509 : std_logic_vector(7 downto 0);
    signal call_225 : std_logic_vector(7 downto 0);
    signal cmp180_738 : std_logic_vector(0 downto 0);
    signal cmp196_788 : std_logic_vector(0 downto 0);
    signal cmp210_839 : std_logic_vector(0 downto 0);
    signal cmp258_1048 : std_logic_vector(0 downto 0);
    signal cmp258x_xnot_1058 : std_logic_vector(0 downto 0);
    signal cmp267_1072 : std_logic_vector(0 downto 0);
    signal cmp274_1118 : std_logic_vector(0 downto 0);
    signal cmp274x_xnot_1128 : std_logic_vector(0 downto 0);
    signal cmp284_1142 : std_logic_vector(0 downto 0);
    signal cmp390_432 : std_logic_vector(0 downto 0);
    signal conv103_531 : std_logic_vector(63 downto 0);
    signal conv109_549 : std_logic_vector(63 downto 0);
    signal conv115_567 : std_logic_vector(63 downto 0);
    signal conv121_585 : std_logic_vector(63 downto 0);
    signal conv127_603 : std_logic_vector(63 downto 0);
    signal conv134_1340 : std_logic_vector(63 downto 0);
    signal conv177_728 : std_logic_vector(31 downto 0);
    signal conv179_646 : std_logic_vector(31 downto 0);
    signal conv189_779 : std_logic_vector(31 downto 0);
    signal conv191_650 : std_logic_vector(31 downto 0);
    signal conv193_654 : std_logic_vector(31 downto 0);
    signal conv19_242 : std_logic_vector(15 downto 0);
    signal conv203_830 : std_logic_vector(31 downto 0);
    signal conv205_669 : std_logic_vector(31 downto 0);
    signal conv22_255 : std_logic_vector(15 downto 0);
    signal conv240_678 : std_logic_vector(15 downto 0);
    signal conv255_1039 : std_logic_vector(31 downto 0);
    signal conv271_1109 : std_logic_vector(31 downto 0);
    signal conv288_1185 : std_logic_vector(31 downto 0);
    signal conv28_267 : std_logic_vector(15 downto 0);
    signal conv294_1232 : std_logic_vector(31 downto 0);
    signal conv300_1278 : std_logic_vector(31 downto 0);
    signal conv310_1348 : std_logic_vector(63 downto 0);
    signal conv317_1357 : std_logic_vector(7 downto 0);
    signal conv31_280 : std_logic_vector(15 downto 0);
    signal conv323_1367 : std_logic_vector(7 downto 0);
    signal conv329_1377 : std_logic_vector(7 downto 0);
    signal conv335_1387 : std_logic_vector(7 downto 0);
    signal conv341_1397 : std_logic_vector(7 downto 0);
    signal conv347_1407 : std_logic_vector(7 downto 0);
    signal conv353_1417 : std_logic_vector(7 downto 0);
    signal conv359_1427 : std_logic_vector(7 downto 0);
    signal conv37_292 : std_logic_vector(15 downto 0);
    signal conv380_1456 : std_logic_vector(31 downto 0);
    signal conv383_1460 : std_logic_vector(31 downto 0);
    signal conv40_305 : std_logic_vector(15 downto 0);
    signal conv47_320 : std_logic_vector(31 downto 0);
    signal conv50_333 : std_logic_vector(31 downto 0);
    signal conv56_345 : std_logic_vector(15 downto 0);
    signal conv59_358 : std_logic_vector(15 downto 0);
    signal conv65_370 : std_logic_vector(15 downto 0);
    signal conv68_383 : std_logic_vector(15 downto 0);
    signal conv73_392 : std_logic_vector(63 downto 0);
    signal conv75_396 : std_logic_vector(63 downto 0);
    signal conv77_400 : std_logic_vector(63 downto 0);
    signal conv79_426 : std_logic_vector(63 downto 0);
    signal conv86_482 : std_logic_vector(63 downto 0);
    signal conv91_495 : std_logic_vector(63 downto 0);
    signal conv97_513 : std_logic_vector(63 downto 0);
    signal exitcond3_623 : std_logic_vector(0 downto 0);
    signal flagx_x0_974 : std_logic_vector(15 downto 0);
    signal i138x_x1_924 : std_logic_vector(15 downto 0);
    signal i138x_x2_714 : std_logic_vector(15 downto 0);
    signal i138x_x2_785_delayed_3_0_802 : std_logic_vector(15 downto 0);
    signal i138x_x2_at_entry_696 : std_logic_vector(15 downto 0);
    signal idxprom290_1207 : std_logic_vector(63 downto 0);
    signal idxprom296_1254 : std_logic_vector(63 downto 0);
    signal idxprom302_1300 : std_logic_vector(63 downto 0);
    signal ifx_xelse292_exec_guard_1098_delayed_1_0_1235 : std_logic_vector(0 downto 0);
    signal ifx_xelse292_exec_guard_1108_delayed_1_0_1248 : std_logic_vector(0 downto 0);
    signal ifx_xelse292_exec_guard_1121_delayed_8_0_1264 : std_logic_vector(0 downto 0);
    signal ifx_xelse292_exec_guard_1132_delayed_1_0_1281 : std_logic_vector(0 downto 0);
    signal ifx_xelse292_exec_guard_1142_delayed_1_0_1294 : std_logic_vector(0 downto 0);
    signal ifx_xelse292_exec_guard_1155_delayed_14_0_1310 : std_logic_vector(0 downto 0);
    signal ifx_xelse292_exec_guard_1223 : std_logic_vector(0 downto 0);
    signal ifx_xelse_exec_guard_764 : std_logic_vector(0 downto 0);
    signal ifx_xelse_exec_guard_771_delayed_1_0_782 : std_logic_vector(0 downto 0);
    signal ifx_xelse_exec_guard_777_delayed_1_0_791 : std_logic_vector(0 downto 0);
    signal ifx_xelse_exec_guard_782_delayed_2_0_799 : std_logic_vector(0 downto 0);
    signal ifx_xelse_exec_guard_788_delayed_1_0_811 : std_logic_vector(0 downto 0);
    signal ifx_xelse_exec_guard_796_delayed_2_0_825 : std_logic_vector(0 downto 0);
    signal ifx_xelse_exec_guard_801_delayed_3_0_833 : std_logic_vector(0 downto 0);
    signal ifx_xelse_exec_guard_808_delayed_3_0_842 : std_logic_vector(0 downto 0);
    signal ifx_xelse_exec_guard_813_delayed_3_0_850 : std_logic_vector(0 downto 0);
    signal ifx_xelse_ifx_xend214_taken_856 : std_logic_vector(0 downto 0);
    signal ifx_xelse_ifx_xthen212_taken_847 : std_logic_vector(0 downto 0);
    signal ifx_xend214_exec_guard_872 : std_logic_vector(0 downto 0);
    signal ifx_xend214_exec_guard_965_delayed_1_0_1042 : std_logic_vector(0 downto 0);
    signal ifx_xend214_exec_guard_971_delayed_1_0_1051 : std_logic_vector(0 downto 0);
    signal ifx_xend214_exec_guard_978_delayed_1_0_1061 : std_logic_vector(0 downto 0);
    signal ifx_xend214_exec_guard_986_delayed_1_0_1075 : std_logic_vector(0 downto 0);
    signal ifx_xend214_exec_guard_993_delayed_1_0_1084 : std_logic_vector(0 downto 0);
    signal ifx_xend214_exec_guard_998_delayed_1_0_1092 : std_logic_vector(0 downto 0);
    signal ifx_xend214_ifx_xthen286_taken_1050_delayed_1_0_1171 : std_logic_vector(0 downto 0);
    signal ifx_xend214_ifx_xthen286_taken_1098 : std_logic_vector(0 downto 0);
    signal ifx_xend214_lorx_xlhsx_xfalse269_taken_1089 : std_logic_vector(0 downto 0);
    signal ifx_xend304_whilex_xend_taken_1328 : std_logic_vector(0 downto 0);
    signal ifx_xthen212_exec_guard_859 : std_logic_vector(0 downto 0);
    signal ifx_xthen212_ifx_xend214_taken_862 : std_logic_vector(0 downto 0);
    signal ifx_xthen286_exec_guard_1060_delayed_1_0_1188 : std_logic_vector(0 downto 0);
    signal ifx_xthen286_exec_guard_1070_delayed_1_0_1201 : std_logic_vector(0 downto 0);
    signal ifx_xthen286_exec_guard_1176 : std_logic_vector(0 downto 0);
    signal ifx_xthen_exec_guard_748 : std_logic_vector(0 downto 0);
    signal ifx_xthen_ifx_xend214_taken_761 : std_logic_vector(0 downto 0);
    signal ifx_xthen_ifx_xend214_taken_826_delayed_3_0_865 : std_logic_vector(0 downto 0);
    signal ifx_xthen_ifx_xend214_taken_832_delayed_3_0_875 : std_logic_vector(0 downto 0);
    signal ifx_xthen_ifx_xend214_taken_850_delayed_3_0_899 : std_logic_vector(0 downto 0);
    signal ifx_xthen_ifx_xend214_taken_866_delayed_3_0_927 : std_logic_vector(0 downto 0);
    signal ifx_xthen_ifx_xend214_taken_882_delayed_3_0_955 : std_logic_vector(0 downto 0);
    signal inc187_774 : std_logic_vector(15 downto 0);
    signal inc187_793_delayed_1_0_814 : std_logic_vector(15 downto 0);
    signal inc201_796 : std_logic_vector(15 downto 0);
    signal inc201x_xi138x_x2_808 : std_logic_vector(15 downto 0);
    signal indvar_461 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_618 : std_logic_vector(63 downto 0);
    signal jx_x0_1008_delayed_1_0_1104 : std_logic_vector(15 downto 0);
    signal jx_x0_952 : std_logic_vector(15 downto 0);
    signal jx_x1_719 : std_logic_vector(15 downto 0);
    signal jx_x1_761_delayed_1_0_767 : std_logic_vector(15 downto 0);
    signal jx_x1_at_entry_701 : std_logic_vector(15 downto 0);
    signal jx_x2_822 : std_logic_vector(15 downto 0);
    signal kx_x0_896 : std_logic_vector(15 downto 0);
    signal kx_x1_709 : std_logic_vector(15 downto 0);
    signal kx_x1_748_delayed_1_0_751 : std_logic_vector(15 downto 0);
    signal kx_x1_at_entry_691 : std_logic_vector(15 downto 0);
    signal lorx_xlhsx_xfalse269_exec_guard_1011_delayed_1_0_1112 : std_logic_vector(0 downto 0);
    signal lorx_xlhsx_xfalse269_exec_guard_1017_delayed_1_0_1121 : std_logic_vector(0 downto 0);
    signal lorx_xlhsx_xfalse269_exec_guard_1024_delayed_1_0_1131 : std_logic_vector(0 downto 0);
    signal lorx_xlhsx_xfalse269_exec_guard_1032_delayed_1_0_1145 : std_logic_vector(0 downto 0);
    signal lorx_xlhsx_xfalse269_exec_guard_1039_delayed_1_0_1154 : std_logic_vector(0 downto 0);
    signal lorx_xlhsx_xfalse269_exec_guard_1044_delayed_1_0_1162 : std_logic_vector(0 downto 0);
    signal lorx_xlhsx_xfalse269_exec_guard_1101 : std_logic_vector(0 downto 0);
    signal lorx_xlhsx_xfalse269_ifx_xelse292_taken_1159 : std_logic_vector(0 downto 0);
    signal lorx_xlhsx_xfalse269_ifx_xthen286_taken_1168 : std_logic_vector(0 downto 0);
    signal mul229_980 : std_logic_vector(15 downto 0);
    signal mul251_1016 : std_logic_vector(15 downto 0);
    signal mul381_1465 : std_logic_vector(31 downto 0);
    signal mul384_1470 : std_logic_vector(31 downto 0);
    signal mul78_411 : std_logic_vector(63 downto 0);
    signal mul_406 : std_logic_vector(63 downto 0);
    signal orx_xcond393_1151 : std_logic_vector(0 downto 0);
    signal orx_xcond_1081 : std_logic_vector(0 downto 0);
    signal ptr_deref_1217_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1217_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1217_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1217_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1217_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1217_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1268_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1268_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1268_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1268_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1268_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1316_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1316_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1316_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1316_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1316_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1316_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_610_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_610_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_610_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_610_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_610_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_610_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext_416 : std_logic_vector(63 downto 0);
    signal shl100_524 : std_logic_vector(63 downto 0);
    signal shl106_542 : std_logic_vector(63 downto 0);
    signal shl112_560 : std_logic_vector(63 downto 0);
    signal shl118_578 : std_logic_vector(63 downto 0);
    signal shl124_596 : std_logic_vector(63 downto 0);
    signal shl194_660 : std_logic_vector(31 downto 0);
    signal shl20_248 : std_logic_vector(15 downto 0);
    signal shl29_273 : std_logic_vector(15 downto 0);
    signal shl38_298 : std_logic_vector(15 downto 0);
    signal shl48_326 : std_logic_vector(31 downto 0);
    signal shl57_351 : std_logic_vector(15 downto 0);
    signal shl66_376 : std_logic_vector(15 downto 0);
    signal shl88_488 : std_logic_vector(63 downto 0);
    signal shl94_506 : std_logic_vector(63 downto 0);
    signal shr289_1198 : std_logic_vector(31 downto 0);
    signal shr295_1245 : std_logic_vector(31 downto 0);
    signal shr301_1291 : std_logic_vector(31 downto 0);
    signal shr320_1363 : std_logic_vector(63 downto 0);
    signal shr326_1373 : std_logic_vector(63 downto 0);
    signal shr332_1383 : std_logic_vector(63 downto 0);
    signal shr338_1393 : std_logic_vector(63 downto 0);
    signal shr344_1403 : std_logic_vector(63 downto 0);
    signal shr350_1413 : std_logic_vector(63 downto 0);
    signal shr356_1423 : std_logic_vector(63 downto 0);
    signal shr_445 : std_logic_vector(63 downto 0);
    signal sub241_1004 : std_logic_vector(15 downto 0);
    signal sub250_1010 : std_logic_vector(15 downto 0);
    signal sub314_1353 : std_logic_vector(63 downto 0);
    signal sub_641 : std_logic_vector(15 downto 0);
    signal tmp1_451 : std_logic_vector(0 downto 0);
    signal tmp298_1269 : std_logic_vector(63 downto 0);
    signal tmp385_992 : std_logic_vector(15 downto 0);
    signal tmp386_1022 : std_logic_vector(15 downto 0);
    signal tmp387_1028 : std_logic_vector(15 downto 0);
    signal tmp_986 : std_logic_vector(15 downto 0);
    signal tobool_1324 : std_logic_vector(0 downto 0);
    signal type_cast_1029_1029_delayed_1_0_1135 : std_logic_vector(31 downto 0);
    signal type_cast_1056_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1069_wire : std_logic_vector(31 downto 0);
    signal type_cast_1126_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1139_wire : std_logic_vector(31 downto 0);
    signal type_cast_1183_wire : std_logic_vector(31 downto 0);
    signal type_cast_1192_wire : std_logic_vector(31 downto 0);
    signal type_cast_1195_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1205_wire : std_logic_vector(63 downto 0);
    signal type_cast_1219_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1230_wire : std_logic_vector(31 downto 0);
    signal type_cast_1239_wire : std_logic_vector(31 downto 0);
    signal type_cast_1242_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1252_wire : std_logic_vector(63 downto 0);
    signal type_cast_1276_wire : std_logic_vector(31 downto 0);
    signal type_cast_1285_wire : std_logic_vector(31 downto 0);
    signal type_cast_1288_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1298_wire : std_logic_vector(63 downto 0);
    signal type_cast_1322_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1338_wire : std_logic_vector(63 downto 0);
    signal type_cast_1346_wire : std_logic_vector(63 downto 0);
    signal type_cast_1361_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1371_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1381_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1391_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1401_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1411_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1421_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_246_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_271_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_296_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_324_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_349_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_374_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_404_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_420_wire : std_logic_vector(63 downto 0);
    signal type_cast_423_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_430_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_443_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_449_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_456_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_465_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_467_wire : std_logic_vector(63 downto 0);
    signal type_cast_486_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_504_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_522_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_540_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_558_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_576_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_594_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_616_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_639_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_644_wire : std_logic_vector(31 downto 0);
    signal type_cast_658_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_712_wire : std_logic_vector(15 downto 0);
    signal type_cast_717_wire : std_logic_vector(15 downto 0);
    signal type_cast_722_wire : std_logic_vector(15 downto 0);
    signal type_cast_733_733_delayed_2_0_732 : std_logic_vector(31 downto 0);
    signal type_cast_735_wire : std_logic_vector(31 downto 0);
    signal type_cast_756_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_772_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_819_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_834_834_delayed_3_0_879 : std_logic_vector(15 downto 0);
    signal type_cast_852_852_delayed_4_0_903 : std_logic_vector(15 downto 0);
    signal type_cast_855_855_delayed_1_0_907 : std_logic_vector(15 downto 0);
    signal type_cast_858_858_delayed_1_0_911 : std_logic_vector(15 downto 0);
    signal type_cast_868_868_delayed_4_0_931 : std_logic_vector(15 downto 0);
    signal type_cast_871_871_delayed_2_0_935 : std_logic_vector(15 downto 0);
    signal type_cast_874_874_delayed_2_0_939 : std_logic_vector(15 downto 0);
    signal type_cast_886_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_890_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_892_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_920_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_948_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_960_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_964_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_968_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_970_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_983_983_delayed_1_0_1065 : std_logic_vector(31 downto 0);
    signal umax2_458 : std_logic_vector(63 downto 0);
    signal whilex_xbody_ifx_xelse_taken_741 : std_logic_vector(0 downto 0);
    signal whilex_xbody_ifx_xthen_taken_745 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    array_obj_ref_1212_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1212_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1212_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1212_resized_base_address <= "00000000000000";
    array_obj_ref_1259_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1259_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1259_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1259_resized_base_address <= "00000000000000";
    array_obj_ref_1305_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1305_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1305_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1305_resized_base_address <= "00000000000000";
    array_obj_ref_473_constant_part_of_offset <= "00000000000000";
    array_obj_ref_473_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_473_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_473_resized_base_address <= "00000000000000";
    i138x_x2_at_entry_696 <= "0000000000000000";
    jx_x1_at_entry_701 <= "0000000000000000";
    kx_x1_at_entry_691 <= "0000000000000000";
    ptr_deref_1217_word_offset_0 <= "00000000000000";
    ptr_deref_1268_word_offset_0 <= "00000000000000";
    ptr_deref_1316_word_offset_0 <= "00000000000000";
    ptr_deref_610_word_offset_0 <= "00000000000000";
    type_cast_1056_wire_constant <= "1";
    type_cast_1126_wire_constant <= "1";
    type_cast_1195_wire_constant <= "00000000000000000000000000000011";
    type_cast_1219_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1242_wire_constant <= "00000000000000000000000000000011";
    type_cast_1288_wire_constant <= "00000000000000000000000000000011";
    type_cast_1322_wire_constant <= "0000000000000000";
    type_cast_1361_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1371_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1381_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1391_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1401_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1411_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1421_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_246_wire_constant <= "0000000000001000";
    type_cast_271_wire_constant <= "0000000000001000";
    type_cast_296_wire_constant <= "0000000000001000";
    type_cast_324_wire_constant <= "00000000000000000000000000001000";
    type_cast_349_wire_constant <= "0000000000001000";
    type_cast_374_wire_constant <= "0000000000001000";
    type_cast_404_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_423_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_430_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000111";
    type_cast_443_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_449_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_456_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_465_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_486_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_504_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_522_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_540_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_558_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_576_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_594_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_616_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_639_wire_constant <= "1111111111111000";
    type_cast_658_wire_constant <= "00000000000000000000000000000001";
    type_cast_756_wire_constant <= "0000000000001000";
    type_cast_772_wire_constant <= "0000000000000001";
    type_cast_819_wire_constant <= "0000000000000000";
    type_cast_886_wire_constant <= "0000000000000000";
    type_cast_890_wire_constant <= "0000000000000000";
    type_cast_892_wire_constant <= "0000000000000000";
    type_cast_920_wire_constant <= "0000000000000000";
    type_cast_948_wire_constant <= "0000000000000000";
    type_cast_960_wire_constant <= "0000000000000000";
    type_cast_964_wire_constant <= "0000000000000001";
    type_cast_968_wire_constant <= "0000000000000000";
    type_cast_970_wire_constant <= "0000000000000000";
    phi_stmt_461: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_465_wire_constant & type_cast_467_wire;
      req <= phi_stmt_461_req_0 & phi_stmt_461_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_461",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_461_ack_0,
          idata => idata,
          odata => indvar_461,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_461
    phi_stmt_709: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_712_wire & kx_x1_at_entry_691;
      req <= phi_stmt_709_req_0 & phi_stmt_709_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_709",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_709_ack_0,
          idata => idata,
          odata => kx_x1_709,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_709
    phi_stmt_714: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_717_wire & i138x_x2_at_entry_696;
      req <= phi_stmt_714_req_0 & phi_stmt_714_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_714",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_714_ack_0,
          idata => idata,
          odata => i138x_x2_714,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_714
    phi_stmt_719: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_722_wire & jx_x1_at_entry_701;
      req <= phi_stmt_719_req_0 & phi_stmt_719_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_719",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_719_ack_0,
          idata => idata,
          odata => jx_x1_719,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_719
    -- flow-through select operator MUX_457_inst
    umax2_458 <= shr_445 when (tmp1_451(0) /=  '0') else type_cast_456_wire_constant;
    -- flow-through select operator MUX_821_inst
    jx_x2_822 <= type_cast_819_wire_constant when (cmp196_788(0) /=  '0') else inc187_793_delayed_1_0_814;
    -- flow-through select operator MUX_893_inst
    MUX_893_wire <= type_cast_890_wire_constant when (ifx_xelse_ifx_xend214_taken_856(0) /=  '0') else type_cast_892_wire_constant;
    -- flow-through select operator MUX_894_inst
    MUX_894_wire <= type_cast_886_wire_constant when (ifx_xthen212_ifx_xend214_taken_862(0) /=  '0') else MUX_893_wire;
    -- flow-through select operator MUX_895_inst
    kx_x0_896 <= type_cast_834_834_delayed_3_0_879 when (ifx_xthen_ifx_xend214_taken_832_delayed_3_0_875(0) /=  '0') else MUX_894_wire;
    -- flow-through select operator MUX_921_inst
    MUX_921_wire <= type_cast_858_858_delayed_1_0_911 when (ifx_xelse_ifx_xend214_taken_856(0) /=  '0') else type_cast_920_wire_constant;
    -- flow-through select operator MUX_922_inst
    MUX_922_wire <= type_cast_855_855_delayed_1_0_907 when (ifx_xthen212_ifx_xend214_taken_862(0) /=  '0') else MUX_921_wire;
    -- flow-through select operator MUX_923_inst
    i138x_x1_924 <= type_cast_852_852_delayed_4_0_903 when (ifx_xthen_ifx_xend214_taken_850_delayed_3_0_899(0) /=  '0') else MUX_922_wire;
    -- flow-through select operator MUX_949_inst
    MUX_949_wire <= type_cast_874_874_delayed_2_0_939 when (ifx_xelse_ifx_xend214_taken_856(0) /=  '0') else type_cast_948_wire_constant;
    -- flow-through select operator MUX_950_inst
    MUX_950_wire <= type_cast_871_871_delayed_2_0_935 when (ifx_xthen212_ifx_xend214_taken_862(0) /=  '0') else MUX_949_wire;
    -- flow-through select operator MUX_951_inst
    jx_x0_952 <= type_cast_868_868_delayed_4_0_931 when (ifx_xthen_ifx_xend214_taken_866_delayed_3_0_927(0) /=  '0') else MUX_950_wire;
    -- flow-through select operator MUX_971_inst
    MUX_971_wire <= type_cast_968_wire_constant when (ifx_xelse_ifx_xend214_taken_856(0) /=  '0') else type_cast_970_wire_constant;
    -- flow-through select operator MUX_972_inst
    MUX_972_wire <= type_cast_964_wire_constant when (ifx_xthen212_ifx_xend214_taken_862(0) /=  '0') else MUX_971_wire;
    -- flow-through select operator MUX_973_inst
    flagx_x0_974 <= type_cast_960_wire_constant when (ifx_xthen_ifx_xend214_taken_882_delayed_3_0_955(0) /=  '0') else MUX_972_wire;
    W_add230_1056_delayed_2_0_1177_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_add230_1056_delayed_2_0_1177_inst_req_0;
      W_add230_1056_delayed_2_0_1177_inst_ack_0<= wack(0);
      rreq(0) <= W_add230_1056_delayed_2_0_1177_inst_req_1;
      W_add230_1056_delayed_2_0_1177_inst_ack_1<= rack(0);
      W_add230_1056_delayed_2_0_1177_inst : InterlockBuffer generic map ( -- 
        name => "W_add230_1056_delayed_2_0_1177_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add230_998,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add230_1056_delayed_2_0_1179,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_add230_1128_delayed_2_0_1270_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_add230_1128_delayed_2_0_1270_inst_req_0;
      W_add230_1128_delayed_2_0_1270_inst_ack_0<= wack(0);
      rreq(0) <= W_add230_1128_delayed_2_0_1270_inst_req_1;
      W_add230_1128_delayed_2_0_1270_inst_ack_1<= rack(0);
      W_add230_1128_delayed_2_0_1270_inst : InterlockBuffer generic map ( -- 
        name => "W_add230_1128_delayed_2_0_1270_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add230_998,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add230_1128_delayed_2_0_1272,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_add252_1094_delayed_2_0_1224_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_add252_1094_delayed_2_0_1224_inst_req_0;
      W_add252_1094_delayed_2_0_1224_inst_ack_0<= wack(0);
      rreq(0) <= W_add252_1094_delayed_2_0_1224_inst_req_1;
      W_add252_1094_delayed_2_0_1224_inst_ack_1<= rack(0);
      W_add252_1094_delayed_2_0_1224_inst : InterlockBuffer generic map ( -- 
        name => "W_add252_1094_delayed_2_0_1224_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add252_1034,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add252_1094_delayed_2_0_1226,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_arrayidx303_1156_delayed_5_0_1311_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_arrayidx303_1156_delayed_5_0_1311_inst_req_0;
      W_arrayidx303_1156_delayed_5_0_1311_inst_ack_0<= wack(0);
      rreq(0) <= W_arrayidx303_1156_delayed_5_0_1311_inst_req_1;
      W_arrayidx303_1156_delayed_5_0_1311_inst_ack_1<= rack(0);
      W_arrayidx303_1156_delayed_5_0_1311_inst : InterlockBuffer generic map ( -- 
        name => "W_arrayidx303_1156_delayed_5_0_1311_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => arrayidx303_1307,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx303_1156_delayed_5_0_1313,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_i138x_x2_785_delayed_3_0_800_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_i138x_x2_785_delayed_3_0_800_inst_req_0;
      W_i138x_x2_785_delayed_3_0_800_inst_ack_0<= wack(0);
      rreq(0) <= W_i138x_x2_785_delayed_3_0_800_inst_req_1;
      W_i138x_x2_785_delayed_3_0_800_inst_ack_1<= rack(0);
      W_i138x_x2_785_delayed_3_0_800_inst : InterlockBuffer generic map ( -- 
        name => "W_i138x_x2_785_delayed_3_0_800_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i138x_x2_714,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => i138x_x2_785_delayed_3_0_802,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xelse292_exec_guard_1098_delayed_1_0_1233_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xelse292_exec_guard_1098_delayed_1_0_1233_inst_req_0;
      W_ifx_xelse292_exec_guard_1098_delayed_1_0_1233_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xelse292_exec_guard_1098_delayed_1_0_1233_inst_req_1;
      W_ifx_xelse292_exec_guard_1098_delayed_1_0_1233_inst_ack_1<= rack(0);
      W_ifx_xelse292_exec_guard_1098_delayed_1_0_1233_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xelse292_exec_guard_1098_delayed_1_0_1233_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xelse292_exec_guard_1223,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xelse292_exec_guard_1098_delayed_1_0_1235,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xelse292_exec_guard_1108_delayed_1_0_1246_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xelse292_exec_guard_1108_delayed_1_0_1246_inst_req_0;
      W_ifx_xelse292_exec_guard_1108_delayed_1_0_1246_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xelse292_exec_guard_1108_delayed_1_0_1246_inst_req_1;
      W_ifx_xelse292_exec_guard_1108_delayed_1_0_1246_inst_ack_1<= rack(0);
      W_ifx_xelse292_exec_guard_1108_delayed_1_0_1246_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xelse292_exec_guard_1108_delayed_1_0_1246_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xelse292_exec_guard_1223,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xelse292_exec_guard_1108_delayed_1_0_1248,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xelse292_exec_guard_1121_delayed_8_0_1262_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xelse292_exec_guard_1121_delayed_8_0_1262_inst_req_0;
      W_ifx_xelse292_exec_guard_1121_delayed_8_0_1262_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xelse292_exec_guard_1121_delayed_8_0_1262_inst_req_1;
      W_ifx_xelse292_exec_guard_1121_delayed_8_0_1262_inst_ack_1<= rack(0);
      W_ifx_xelse292_exec_guard_1121_delayed_8_0_1262_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xelse292_exec_guard_1121_delayed_8_0_1262_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xelse292_exec_guard_1223,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xelse292_exec_guard_1121_delayed_8_0_1264,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xelse292_exec_guard_1132_delayed_1_0_1279_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xelse292_exec_guard_1132_delayed_1_0_1279_inst_req_0;
      W_ifx_xelse292_exec_guard_1132_delayed_1_0_1279_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xelse292_exec_guard_1132_delayed_1_0_1279_inst_req_1;
      W_ifx_xelse292_exec_guard_1132_delayed_1_0_1279_inst_ack_1<= rack(0);
      W_ifx_xelse292_exec_guard_1132_delayed_1_0_1279_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xelse292_exec_guard_1132_delayed_1_0_1279_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xelse292_exec_guard_1223,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xelse292_exec_guard_1132_delayed_1_0_1281,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xelse292_exec_guard_1142_delayed_1_0_1292_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xelse292_exec_guard_1142_delayed_1_0_1292_inst_req_0;
      W_ifx_xelse292_exec_guard_1142_delayed_1_0_1292_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xelse292_exec_guard_1142_delayed_1_0_1292_inst_req_1;
      W_ifx_xelse292_exec_guard_1142_delayed_1_0_1292_inst_ack_1<= rack(0);
      W_ifx_xelse292_exec_guard_1142_delayed_1_0_1292_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xelse292_exec_guard_1142_delayed_1_0_1292_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xelse292_exec_guard_1223,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xelse292_exec_guard_1142_delayed_1_0_1294,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xelse292_exec_guard_1155_delayed_14_0_1308_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xelse292_exec_guard_1155_delayed_14_0_1308_inst_req_0;
      W_ifx_xelse292_exec_guard_1155_delayed_14_0_1308_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xelse292_exec_guard_1155_delayed_14_0_1308_inst_req_1;
      W_ifx_xelse292_exec_guard_1155_delayed_14_0_1308_inst_ack_1<= rack(0);
      W_ifx_xelse292_exec_guard_1155_delayed_14_0_1308_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xelse292_exec_guard_1155_delayed_14_0_1308_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xelse292_exec_guard_1223,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xelse292_exec_guard_1155_delayed_14_0_1310,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_ifx_xelse292_exec_guard_1221_inst
    process(lorx_xlhsx_xfalse269_ifx_xelse292_taken_1159) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := lorx_xlhsx_xfalse269_ifx_xelse292_taken_1159(0 downto 0);
      ifx_xelse292_exec_guard_1223 <= tmp_var; -- 
    end process;
    -- interlock W_ifx_xelse_exec_guard_762_inst
    process(whilex_xbody_ifx_xelse_taken_741) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := whilex_xbody_ifx_xelse_taken_741(0 downto 0);
      ifx_xelse_exec_guard_764 <= tmp_var; -- 
    end process;
    W_ifx_xelse_exec_guard_771_delayed_1_0_780_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xelse_exec_guard_771_delayed_1_0_780_inst_req_0;
      W_ifx_xelse_exec_guard_771_delayed_1_0_780_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xelse_exec_guard_771_delayed_1_0_780_inst_req_1;
      W_ifx_xelse_exec_guard_771_delayed_1_0_780_inst_ack_1<= rack(0);
      W_ifx_xelse_exec_guard_771_delayed_1_0_780_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xelse_exec_guard_771_delayed_1_0_780_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xelse_exec_guard_764,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xelse_exec_guard_771_delayed_1_0_782,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xelse_exec_guard_777_delayed_1_0_789_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xelse_exec_guard_777_delayed_1_0_789_inst_req_0;
      W_ifx_xelse_exec_guard_777_delayed_1_0_789_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xelse_exec_guard_777_delayed_1_0_789_inst_req_1;
      W_ifx_xelse_exec_guard_777_delayed_1_0_789_inst_ack_1<= rack(0);
      W_ifx_xelse_exec_guard_777_delayed_1_0_789_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xelse_exec_guard_777_delayed_1_0_789_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xelse_exec_guard_764,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xelse_exec_guard_777_delayed_1_0_791,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xelse_exec_guard_782_delayed_2_0_797_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xelse_exec_guard_782_delayed_2_0_797_inst_req_0;
      W_ifx_xelse_exec_guard_782_delayed_2_0_797_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xelse_exec_guard_782_delayed_2_0_797_inst_req_1;
      W_ifx_xelse_exec_guard_782_delayed_2_0_797_inst_ack_1<= rack(0);
      W_ifx_xelse_exec_guard_782_delayed_2_0_797_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xelse_exec_guard_782_delayed_2_0_797_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xelse_exec_guard_764,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xelse_exec_guard_782_delayed_2_0_799,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xelse_exec_guard_788_delayed_1_0_809_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xelse_exec_guard_788_delayed_1_0_809_inst_req_0;
      W_ifx_xelse_exec_guard_788_delayed_1_0_809_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xelse_exec_guard_788_delayed_1_0_809_inst_req_1;
      W_ifx_xelse_exec_guard_788_delayed_1_0_809_inst_ack_1<= rack(0);
      W_ifx_xelse_exec_guard_788_delayed_1_0_809_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xelse_exec_guard_788_delayed_1_0_809_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xelse_exec_guard_764,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xelse_exec_guard_788_delayed_1_0_811,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xelse_exec_guard_796_delayed_2_0_823_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xelse_exec_guard_796_delayed_2_0_823_inst_req_0;
      W_ifx_xelse_exec_guard_796_delayed_2_0_823_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xelse_exec_guard_796_delayed_2_0_823_inst_req_1;
      W_ifx_xelse_exec_guard_796_delayed_2_0_823_inst_ack_1<= rack(0);
      W_ifx_xelse_exec_guard_796_delayed_2_0_823_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xelse_exec_guard_796_delayed_2_0_823_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xelse_exec_guard_764,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xelse_exec_guard_796_delayed_2_0_825,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xelse_exec_guard_801_delayed_3_0_831_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xelse_exec_guard_801_delayed_3_0_831_inst_req_0;
      W_ifx_xelse_exec_guard_801_delayed_3_0_831_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xelse_exec_guard_801_delayed_3_0_831_inst_req_1;
      W_ifx_xelse_exec_guard_801_delayed_3_0_831_inst_ack_1<= rack(0);
      W_ifx_xelse_exec_guard_801_delayed_3_0_831_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xelse_exec_guard_801_delayed_3_0_831_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xelse_exec_guard_764,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xelse_exec_guard_801_delayed_3_0_833,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xelse_exec_guard_808_delayed_3_0_840_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xelse_exec_guard_808_delayed_3_0_840_inst_req_0;
      W_ifx_xelse_exec_guard_808_delayed_3_0_840_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xelse_exec_guard_808_delayed_3_0_840_inst_req_1;
      W_ifx_xelse_exec_guard_808_delayed_3_0_840_inst_ack_1<= rack(0);
      W_ifx_xelse_exec_guard_808_delayed_3_0_840_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xelse_exec_guard_808_delayed_3_0_840_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xelse_exec_guard_764,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xelse_exec_guard_808_delayed_3_0_842,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xelse_exec_guard_813_delayed_3_0_848_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xelse_exec_guard_813_delayed_3_0_848_inst_req_0;
      W_ifx_xelse_exec_guard_813_delayed_3_0_848_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xelse_exec_guard_813_delayed_3_0_848_inst_req_1;
      W_ifx_xelse_exec_guard_813_delayed_3_0_848_inst_ack_1<= rack(0);
      W_ifx_xelse_exec_guard_813_delayed_3_0_848_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xelse_exec_guard_813_delayed_3_0_848_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xelse_exec_guard_764,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xelse_exec_guard_813_delayed_3_0_850,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xend214_exec_guard_965_delayed_1_0_1040_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xend214_exec_guard_965_delayed_1_0_1040_inst_req_0;
      W_ifx_xend214_exec_guard_965_delayed_1_0_1040_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xend214_exec_guard_965_delayed_1_0_1040_inst_req_1;
      W_ifx_xend214_exec_guard_965_delayed_1_0_1040_inst_ack_1<= rack(0);
      W_ifx_xend214_exec_guard_965_delayed_1_0_1040_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xend214_exec_guard_965_delayed_1_0_1040_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xend214_exec_guard_872,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xend214_exec_guard_965_delayed_1_0_1042,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xend214_exec_guard_971_delayed_1_0_1049_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xend214_exec_guard_971_delayed_1_0_1049_inst_req_0;
      W_ifx_xend214_exec_guard_971_delayed_1_0_1049_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xend214_exec_guard_971_delayed_1_0_1049_inst_req_1;
      W_ifx_xend214_exec_guard_971_delayed_1_0_1049_inst_ack_1<= rack(0);
      W_ifx_xend214_exec_guard_971_delayed_1_0_1049_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xend214_exec_guard_971_delayed_1_0_1049_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xend214_exec_guard_872,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xend214_exec_guard_971_delayed_1_0_1051,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xend214_exec_guard_978_delayed_1_0_1059_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xend214_exec_guard_978_delayed_1_0_1059_inst_req_0;
      W_ifx_xend214_exec_guard_978_delayed_1_0_1059_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xend214_exec_guard_978_delayed_1_0_1059_inst_req_1;
      W_ifx_xend214_exec_guard_978_delayed_1_0_1059_inst_ack_1<= rack(0);
      W_ifx_xend214_exec_guard_978_delayed_1_0_1059_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xend214_exec_guard_978_delayed_1_0_1059_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xend214_exec_guard_872,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xend214_exec_guard_978_delayed_1_0_1061,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xend214_exec_guard_986_delayed_1_0_1073_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xend214_exec_guard_986_delayed_1_0_1073_inst_req_0;
      W_ifx_xend214_exec_guard_986_delayed_1_0_1073_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xend214_exec_guard_986_delayed_1_0_1073_inst_req_1;
      W_ifx_xend214_exec_guard_986_delayed_1_0_1073_inst_ack_1<= rack(0);
      W_ifx_xend214_exec_guard_986_delayed_1_0_1073_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xend214_exec_guard_986_delayed_1_0_1073_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xend214_exec_guard_872,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xend214_exec_guard_986_delayed_1_0_1075,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xend214_exec_guard_993_delayed_1_0_1082_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xend214_exec_guard_993_delayed_1_0_1082_inst_req_0;
      W_ifx_xend214_exec_guard_993_delayed_1_0_1082_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xend214_exec_guard_993_delayed_1_0_1082_inst_req_1;
      W_ifx_xend214_exec_guard_993_delayed_1_0_1082_inst_ack_1<= rack(0);
      W_ifx_xend214_exec_guard_993_delayed_1_0_1082_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xend214_exec_guard_993_delayed_1_0_1082_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xend214_exec_guard_872,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xend214_exec_guard_993_delayed_1_0_1084,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xend214_exec_guard_998_delayed_1_0_1090_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xend214_exec_guard_998_delayed_1_0_1090_inst_req_0;
      W_ifx_xend214_exec_guard_998_delayed_1_0_1090_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xend214_exec_guard_998_delayed_1_0_1090_inst_req_1;
      W_ifx_xend214_exec_guard_998_delayed_1_0_1090_inst_ack_1<= rack(0);
      W_ifx_xend214_exec_guard_998_delayed_1_0_1090_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xend214_exec_guard_998_delayed_1_0_1090_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xend214_exec_guard_872,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xend214_exec_guard_998_delayed_1_0_1092,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xend214_ifx_xthen286_taken_1050_delayed_1_0_1169_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xend214_ifx_xthen286_taken_1050_delayed_1_0_1169_inst_req_0;
      W_ifx_xend214_ifx_xthen286_taken_1050_delayed_1_0_1169_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xend214_ifx_xthen286_taken_1050_delayed_1_0_1169_inst_req_1;
      W_ifx_xend214_ifx_xthen286_taken_1050_delayed_1_0_1169_inst_ack_1<= rack(0);
      W_ifx_xend214_ifx_xthen286_taken_1050_delayed_1_0_1169_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xend214_ifx_xthen286_taken_1050_delayed_1_0_1169_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xend214_ifx_xthen286_taken_1098,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xend214_ifx_xthen286_taken_1050_delayed_1_0_1171,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_ifx_xthen212_exec_guard_857_inst
    process(ifx_xelse_ifx_xthen212_taken_847) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := ifx_xelse_ifx_xthen212_taken_847(0 downto 0);
      ifx_xthen212_exec_guard_859 <= tmp_var; -- 
    end process;
    -- interlock W_ifx_xthen212_ifx_xend214_taken_860_inst
    process(ifx_xthen212_exec_guard_859) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := ifx_xthen212_exec_guard_859(0 downto 0);
      ifx_xthen212_ifx_xend214_taken_862 <= tmp_var; -- 
    end process;
    W_ifx_xthen286_exec_guard_1060_delayed_1_0_1186_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xthen286_exec_guard_1060_delayed_1_0_1186_inst_req_0;
      W_ifx_xthen286_exec_guard_1060_delayed_1_0_1186_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xthen286_exec_guard_1060_delayed_1_0_1186_inst_req_1;
      W_ifx_xthen286_exec_guard_1060_delayed_1_0_1186_inst_ack_1<= rack(0);
      W_ifx_xthen286_exec_guard_1060_delayed_1_0_1186_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xthen286_exec_guard_1060_delayed_1_0_1186_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xthen286_exec_guard_1176,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xthen286_exec_guard_1060_delayed_1_0_1188,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xthen286_exec_guard_1070_delayed_1_0_1199_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xthen286_exec_guard_1070_delayed_1_0_1199_inst_req_0;
      W_ifx_xthen286_exec_guard_1070_delayed_1_0_1199_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xthen286_exec_guard_1070_delayed_1_0_1199_inst_req_1;
      W_ifx_xthen286_exec_guard_1070_delayed_1_0_1199_inst_ack_1<= rack(0);
      W_ifx_xthen286_exec_guard_1070_delayed_1_0_1199_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xthen286_exec_guard_1070_delayed_1_0_1199_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xthen286_exec_guard_1176,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xthen286_exec_guard_1070_delayed_1_0_1201,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_ifx_xthen_exec_guard_746_inst
    process(whilex_xbody_ifx_xthen_taken_745) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := whilex_xbody_ifx_xthen_taken_745(0 downto 0);
      ifx_xthen_exec_guard_748 <= tmp_var; -- 
    end process;
    -- interlock W_ifx_xthen_ifx_xend214_taken_759_inst
    process(ifx_xthen_exec_guard_748) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := ifx_xthen_exec_guard_748(0 downto 0);
      ifx_xthen_ifx_xend214_taken_761 <= tmp_var; -- 
    end process;
    W_ifx_xthen_ifx_xend214_taken_826_delayed_3_0_863_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xthen_ifx_xend214_taken_826_delayed_3_0_863_inst_req_0;
      W_ifx_xthen_ifx_xend214_taken_826_delayed_3_0_863_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xthen_ifx_xend214_taken_826_delayed_3_0_863_inst_req_1;
      W_ifx_xthen_ifx_xend214_taken_826_delayed_3_0_863_inst_ack_1<= rack(0);
      W_ifx_xthen_ifx_xend214_taken_826_delayed_3_0_863_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xthen_ifx_xend214_taken_826_delayed_3_0_863_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xthen_ifx_xend214_taken_761,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xthen_ifx_xend214_taken_826_delayed_3_0_865,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xthen_ifx_xend214_taken_832_delayed_3_0_873_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xthen_ifx_xend214_taken_832_delayed_3_0_873_inst_req_0;
      W_ifx_xthen_ifx_xend214_taken_832_delayed_3_0_873_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xthen_ifx_xend214_taken_832_delayed_3_0_873_inst_req_1;
      W_ifx_xthen_ifx_xend214_taken_832_delayed_3_0_873_inst_ack_1<= rack(0);
      W_ifx_xthen_ifx_xend214_taken_832_delayed_3_0_873_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xthen_ifx_xend214_taken_832_delayed_3_0_873_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xthen_ifx_xend214_taken_761,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xthen_ifx_xend214_taken_832_delayed_3_0_875,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xthen_ifx_xend214_taken_850_delayed_3_0_897_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xthen_ifx_xend214_taken_850_delayed_3_0_897_inst_req_0;
      W_ifx_xthen_ifx_xend214_taken_850_delayed_3_0_897_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xthen_ifx_xend214_taken_850_delayed_3_0_897_inst_req_1;
      W_ifx_xthen_ifx_xend214_taken_850_delayed_3_0_897_inst_ack_1<= rack(0);
      W_ifx_xthen_ifx_xend214_taken_850_delayed_3_0_897_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xthen_ifx_xend214_taken_850_delayed_3_0_897_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xthen_ifx_xend214_taken_761,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xthen_ifx_xend214_taken_850_delayed_3_0_899,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xthen_ifx_xend214_taken_866_delayed_3_0_925_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xthen_ifx_xend214_taken_866_delayed_3_0_925_inst_req_0;
      W_ifx_xthen_ifx_xend214_taken_866_delayed_3_0_925_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xthen_ifx_xend214_taken_866_delayed_3_0_925_inst_req_1;
      W_ifx_xthen_ifx_xend214_taken_866_delayed_3_0_925_inst_ack_1<= rack(0);
      W_ifx_xthen_ifx_xend214_taken_866_delayed_3_0_925_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xthen_ifx_xend214_taken_866_delayed_3_0_925_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xthen_ifx_xend214_taken_761,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xthen_ifx_xend214_taken_866_delayed_3_0_927,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xthen_ifx_xend214_taken_882_delayed_3_0_953_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xthen_ifx_xend214_taken_882_delayed_3_0_953_inst_req_0;
      W_ifx_xthen_ifx_xend214_taken_882_delayed_3_0_953_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xthen_ifx_xend214_taken_882_delayed_3_0_953_inst_req_1;
      W_ifx_xthen_ifx_xend214_taken_882_delayed_3_0_953_inst_ack_1<= rack(0);
      W_ifx_xthen_ifx_xend214_taken_882_delayed_3_0_953_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xthen_ifx_xend214_taken_882_delayed_3_0_953_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xthen_ifx_xend214_taken_761,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xthen_ifx_xend214_taken_882_delayed_3_0_955,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_inc187_793_delayed_1_0_812_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_inc187_793_delayed_1_0_812_inst_req_0;
      W_inc187_793_delayed_1_0_812_inst_ack_0<= wack(0);
      rreq(0) <= W_inc187_793_delayed_1_0_812_inst_req_1;
      W_inc187_793_delayed_1_0_812_inst_ack_1<= rack(0);
      W_inc187_793_delayed_1_0_812_inst : InterlockBuffer generic map ( -- 
        name => "W_inc187_793_delayed_1_0_812_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc187_774,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc187_793_delayed_1_0_814,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_jx_x0_1008_delayed_1_0_1102_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_jx_x0_1008_delayed_1_0_1102_inst_req_0;
      W_jx_x0_1008_delayed_1_0_1102_inst_ack_0<= wack(0);
      rreq(0) <= W_jx_x0_1008_delayed_1_0_1102_inst_req_1;
      W_jx_x0_1008_delayed_1_0_1102_inst_ack_1<= rack(0);
      W_jx_x0_1008_delayed_1_0_1102_inst : InterlockBuffer generic map ( -- 
        name => "W_jx_x0_1008_delayed_1_0_1102_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x0_952,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => jx_x0_1008_delayed_1_0_1104,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_jx_x1_761_delayed_1_0_765_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_jx_x1_761_delayed_1_0_765_inst_req_0;
      W_jx_x1_761_delayed_1_0_765_inst_ack_0<= wack(0);
      rreq(0) <= W_jx_x1_761_delayed_1_0_765_inst_req_1;
      W_jx_x1_761_delayed_1_0_765_inst_ack_1<= rack(0);
      W_jx_x1_761_delayed_1_0_765_inst : InterlockBuffer generic map ( -- 
        name => "W_jx_x1_761_delayed_1_0_765_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x1_719,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => jx_x1_761_delayed_1_0_767,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_kx_x1_748_delayed_1_0_749_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_kx_x1_748_delayed_1_0_749_inst_req_0;
      W_kx_x1_748_delayed_1_0_749_inst_ack_0<= wack(0);
      rreq(0) <= W_kx_x1_748_delayed_1_0_749_inst_req_1;
      W_kx_x1_748_delayed_1_0_749_inst_ack_1<= rack(0);
      W_kx_x1_748_delayed_1_0_749_inst : InterlockBuffer generic map ( -- 
        name => "W_kx_x1_748_delayed_1_0_749_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => kx_x1_709,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => kx_x1_748_delayed_1_0_751,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_lorx_xlhsx_xfalse269_exec_guard_1011_delayed_1_0_1110_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_lorx_xlhsx_xfalse269_exec_guard_1011_delayed_1_0_1110_inst_req_0;
      W_lorx_xlhsx_xfalse269_exec_guard_1011_delayed_1_0_1110_inst_ack_0<= wack(0);
      rreq(0) <= W_lorx_xlhsx_xfalse269_exec_guard_1011_delayed_1_0_1110_inst_req_1;
      W_lorx_xlhsx_xfalse269_exec_guard_1011_delayed_1_0_1110_inst_ack_1<= rack(0);
      W_lorx_xlhsx_xfalse269_exec_guard_1011_delayed_1_0_1110_inst : InterlockBuffer generic map ( -- 
        name => "W_lorx_xlhsx_xfalse269_exec_guard_1011_delayed_1_0_1110_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => lorx_xlhsx_xfalse269_exec_guard_1101,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => lorx_xlhsx_xfalse269_exec_guard_1011_delayed_1_0_1112,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_lorx_xlhsx_xfalse269_exec_guard_1017_delayed_1_0_1119_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_lorx_xlhsx_xfalse269_exec_guard_1017_delayed_1_0_1119_inst_req_0;
      W_lorx_xlhsx_xfalse269_exec_guard_1017_delayed_1_0_1119_inst_ack_0<= wack(0);
      rreq(0) <= W_lorx_xlhsx_xfalse269_exec_guard_1017_delayed_1_0_1119_inst_req_1;
      W_lorx_xlhsx_xfalse269_exec_guard_1017_delayed_1_0_1119_inst_ack_1<= rack(0);
      W_lorx_xlhsx_xfalse269_exec_guard_1017_delayed_1_0_1119_inst : InterlockBuffer generic map ( -- 
        name => "W_lorx_xlhsx_xfalse269_exec_guard_1017_delayed_1_0_1119_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => lorx_xlhsx_xfalse269_exec_guard_1101,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => lorx_xlhsx_xfalse269_exec_guard_1017_delayed_1_0_1121,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_lorx_xlhsx_xfalse269_exec_guard_1024_delayed_1_0_1129_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_lorx_xlhsx_xfalse269_exec_guard_1024_delayed_1_0_1129_inst_req_0;
      W_lorx_xlhsx_xfalse269_exec_guard_1024_delayed_1_0_1129_inst_ack_0<= wack(0);
      rreq(0) <= W_lorx_xlhsx_xfalse269_exec_guard_1024_delayed_1_0_1129_inst_req_1;
      W_lorx_xlhsx_xfalse269_exec_guard_1024_delayed_1_0_1129_inst_ack_1<= rack(0);
      W_lorx_xlhsx_xfalse269_exec_guard_1024_delayed_1_0_1129_inst : InterlockBuffer generic map ( -- 
        name => "W_lorx_xlhsx_xfalse269_exec_guard_1024_delayed_1_0_1129_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => lorx_xlhsx_xfalse269_exec_guard_1101,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => lorx_xlhsx_xfalse269_exec_guard_1024_delayed_1_0_1131,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_lorx_xlhsx_xfalse269_exec_guard_1032_delayed_1_0_1143_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_lorx_xlhsx_xfalse269_exec_guard_1032_delayed_1_0_1143_inst_req_0;
      W_lorx_xlhsx_xfalse269_exec_guard_1032_delayed_1_0_1143_inst_ack_0<= wack(0);
      rreq(0) <= W_lorx_xlhsx_xfalse269_exec_guard_1032_delayed_1_0_1143_inst_req_1;
      W_lorx_xlhsx_xfalse269_exec_guard_1032_delayed_1_0_1143_inst_ack_1<= rack(0);
      W_lorx_xlhsx_xfalse269_exec_guard_1032_delayed_1_0_1143_inst : InterlockBuffer generic map ( -- 
        name => "W_lorx_xlhsx_xfalse269_exec_guard_1032_delayed_1_0_1143_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => lorx_xlhsx_xfalse269_exec_guard_1101,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => lorx_xlhsx_xfalse269_exec_guard_1032_delayed_1_0_1145,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_lorx_xlhsx_xfalse269_exec_guard_1039_delayed_1_0_1152_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_lorx_xlhsx_xfalse269_exec_guard_1039_delayed_1_0_1152_inst_req_0;
      W_lorx_xlhsx_xfalse269_exec_guard_1039_delayed_1_0_1152_inst_ack_0<= wack(0);
      rreq(0) <= W_lorx_xlhsx_xfalse269_exec_guard_1039_delayed_1_0_1152_inst_req_1;
      W_lorx_xlhsx_xfalse269_exec_guard_1039_delayed_1_0_1152_inst_ack_1<= rack(0);
      W_lorx_xlhsx_xfalse269_exec_guard_1039_delayed_1_0_1152_inst : InterlockBuffer generic map ( -- 
        name => "W_lorx_xlhsx_xfalse269_exec_guard_1039_delayed_1_0_1152_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => lorx_xlhsx_xfalse269_exec_guard_1101,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => lorx_xlhsx_xfalse269_exec_guard_1039_delayed_1_0_1154,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_lorx_xlhsx_xfalse269_exec_guard_1044_delayed_1_0_1160_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_lorx_xlhsx_xfalse269_exec_guard_1044_delayed_1_0_1160_inst_req_0;
      W_lorx_xlhsx_xfalse269_exec_guard_1044_delayed_1_0_1160_inst_ack_0<= wack(0);
      rreq(0) <= W_lorx_xlhsx_xfalse269_exec_guard_1044_delayed_1_0_1160_inst_req_1;
      W_lorx_xlhsx_xfalse269_exec_guard_1044_delayed_1_0_1160_inst_ack_1<= rack(0);
      W_lorx_xlhsx_xfalse269_exec_guard_1044_delayed_1_0_1160_inst : InterlockBuffer generic map ( -- 
        name => "W_lorx_xlhsx_xfalse269_exec_guard_1044_delayed_1_0_1160_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => lorx_xlhsx_xfalse269_exec_guard_1101,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => lorx_xlhsx_xfalse269_exec_guard_1044_delayed_1_0_1162,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_lorx_xlhsx_xfalse269_exec_guard_1099_inst
    process(ifx_xend214_lorx_xlhsx_xfalse269_taken_1089) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := ifx_xend214_lorx_xlhsx_xfalse269_taken_1089(0 downto 0);
      lorx_xlhsx_xfalse269_exec_guard_1101 <= tmp_var; -- 
    end process;
    -- interlock W_whilex_xbody_ifx_xelse_taken_739_inst
    process(cmp180_738) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := cmp180_738(0 downto 0);
      whilex_xbody_ifx_xelse_taken_741 <= tmp_var; -- 
    end process;
    addr_of_1213_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1213_final_reg_req_0;
      addr_of_1213_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1213_final_reg_req_1;
      addr_of_1213_final_reg_ack_1<= rack(0);
      addr_of_1213_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1213_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1212_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx291_1214,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1260_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1260_final_reg_req_0;
      addr_of_1260_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1260_final_reg_req_1;
      addr_of_1260_final_reg_ack_1<= rack(0);
      addr_of_1260_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1260_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1259_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx297_1261,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1306_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1306_final_reg_req_0;
      addr_of_1306_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1306_final_reg_req_1;
      addr_of_1306_final_reg_ack_1<= rack(0);
      addr_of_1306_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1306_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1305_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx303_1307,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_474_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_474_final_reg_req_0;
      addr_of_474_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_474_final_reg_req_1;
      addr_of_474_final_reg_ack_1<= rack(0);
      addr_of_474_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_474_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_473_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_475,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1038_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1038_inst_req_0;
      type_cast_1038_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1038_inst_req_1;
      type_cast_1038_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  ifx_xend214_exec_guard_872(0);
      type_cast_1038_inst_gI: SplitGuardInterface generic map(name => "type_cast_1038_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1038_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1038_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i138x_x1_924,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv255_1039,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1064_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1064_inst_req_0;
      type_cast_1064_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1064_inst_req_1;
      type_cast_1064_inst_ack_1<= rack(0);
      type_cast_1064_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1064_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add266_683,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_983_983_delayed_1_0_1065,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1069_inst
    process(conv255_1039) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv255_1039(31 downto 0);
      type_cast_1069_wire <= tmp_var; -- 
    end process;
    type_cast_1108_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1108_inst_req_0;
      type_cast_1108_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1108_inst_req_1;
      type_cast_1108_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  lorx_xlhsx_xfalse269_exec_guard_1101(0);
      type_cast_1108_inst_gI: SplitGuardInterface generic map(name => "type_cast_1108_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1108_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1108_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x0_1008_delayed_1_0_1104,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv271_1109,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1134_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1134_inst_req_0;
      type_cast_1134_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1134_inst_req_1;
      type_cast_1134_inst_ack_1<= rack(0);
      type_cast_1134_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1134_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add283_688,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1029_1029_delayed_1_0_1135,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1139_inst
    process(conv271_1109) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv271_1109(31 downto 0);
      type_cast_1139_wire <= tmp_var; -- 
    end process;
    type_cast_1184_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1184_inst_req_0;
      type_cast_1184_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1184_inst_req_1;
      type_cast_1184_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  ifx_xthen286_exec_guard_1176(0);
      type_cast_1184_inst_gI: SplitGuardInterface generic map(name => "type_cast_1184_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1184_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1184_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1183_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv288_1185,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1192_inst
    process(conv288_1185) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv288_1185(31 downto 0);
      type_cast_1192_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1197_inst
    process(ASHR_i32_i32_1196_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1196_wire(31 downto 0);
      shr289_1198 <= tmp_var; -- 
    end process;
    type_cast_1206_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1206_inst_req_0;
      type_cast_1206_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1206_inst_req_1;
      type_cast_1206_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  ifx_xthen286_exec_guard_1070_delayed_1_0_1201(0);
      type_cast_1206_inst_gI: SplitGuardInterface generic map(name => "type_cast_1206_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1206_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1206_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1205_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom290_1207,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1231_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1231_inst_req_0;
      type_cast_1231_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1231_inst_req_1;
      type_cast_1231_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  ifx_xelse292_exec_guard_1223(0);
      type_cast_1231_inst_gI: SplitGuardInterface generic map(name => "type_cast_1231_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1231_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1231_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1230_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv294_1232,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1239_inst
    process(conv294_1232) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv294_1232(31 downto 0);
      type_cast_1239_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1244_inst
    process(ASHR_i32_i32_1243_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1243_wire(31 downto 0);
      shr295_1245 <= tmp_var; -- 
    end process;
    type_cast_1253_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1253_inst_req_0;
      type_cast_1253_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1253_inst_req_1;
      type_cast_1253_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  ifx_xelse292_exec_guard_1108_delayed_1_0_1248(0);
      type_cast_1253_inst_gI: SplitGuardInterface generic map(name => "type_cast_1253_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1253_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1253_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1252_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom296_1254,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1277_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1277_inst_req_0;
      type_cast_1277_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1277_inst_req_1;
      type_cast_1277_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  ifx_xelse292_exec_guard_1223(0);
      type_cast_1277_inst_gI: SplitGuardInterface generic map(name => "type_cast_1277_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1277_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1277_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1276_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv300_1278,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1285_inst
    process(conv300_1278) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv300_1278(31 downto 0);
      type_cast_1285_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1290_inst
    process(ASHR_i32_i32_1289_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1289_wire(31 downto 0);
      shr301_1291 <= tmp_var; -- 
    end process;
    type_cast_1299_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1299_inst_req_0;
      type_cast_1299_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1299_inst_req_1;
      type_cast_1299_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  ifx_xelse292_exec_guard_1142_delayed_1_0_1294(0);
      type_cast_1299_inst_gI: SplitGuardInterface generic map(name => "type_cast_1299_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1299_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1299_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1298_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom302_1300,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1339_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1339_inst_req_0;
      type_cast_1339_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1339_inst_req_1;
      type_cast_1339_inst_ack_1<= rack(0);
      type_cast_1339_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1339_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1338_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv134_1340,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1347_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1347_inst_req_0;
      type_cast_1347_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1347_inst_req_1;
      type_cast_1347_inst_ack_1<= rack(0);
      type_cast_1347_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1347_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1346_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv310_1348,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1356_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1356_inst_req_0;
      type_cast_1356_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1356_inst_req_1;
      type_cast_1356_inst_ack_1<= rack(0);
      type_cast_1356_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1356_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub314_1353,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv317_1357,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1366_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1366_inst_req_0;
      type_cast_1366_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1366_inst_req_1;
      type_cast_1366_inst_ack_1<= rack(0);
      type_cast_1366_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1366_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr320_1363,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv323_1367,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1376_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1376_inst_req_0;
      type_cast_1376_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1376_inst_req_1;
      type_cast_1376_inst_ack_1<= rack(0);
      type_cast_1376_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1376_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr326_1373,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv329_1377,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1386_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1386_inst_req_0;
      type_cast_1386_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1386_inst_req_1;
      type_cast_1386_inst_ack_1<= rack(0);
      type_cast_1386_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1386_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr332_1383,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv335_1387,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1396_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1396_inst_req_0;
      type_cast_1396_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1396_inst_req_1;
      type_cast_1396_inst_ack_1<= rack(0);
      type_cast_1396_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1396_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr338_1393,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv341_1397,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1406_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1406_inst_req_0;
      type_cast_1406_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1406_inst_req_1;
      type_cast_1406_inst_ack_1<= rack(0);
      type_cast_1406_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1406_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr344_1403,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv347_1407,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1416_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1416_inst_req_0;
      type_cast_1416_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1416_inst_req_1;
      type_cast_1416_inst_ack_1<= rack(0);
      type_cast_1416_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1416_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr350_1413,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv353_1417,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1426_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1426_inst_req_0;
      type_cast_1426_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1426_inst_req_1;
      type_cast_1426_inst_ack_1<= rack(0);
      type_cast_1426_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1426_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr356_1423,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv359_1427,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1455_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1455_inst_req_0;
      type_cast_1455_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1455_inst_req_1;
      type_cast_1455_inst_ack_1<= rack(0);
      type_cast_1455_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1455_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add60_363,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv380_1456,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1459_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1459_inst_req_0;
      type_cast_1459_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1459_inst_req_1;
      type_cast_1459_inst_ack_1<= rack(0);
      type_cast_1459_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1459_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add69_388,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv383_1460,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_241_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_241_inst_req_0;
      type_cast_241_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_241_inst_req_1;
      type_cast_241_inst_ack_1<= rack(0);
      type_cast_241_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_241_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_237,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv19_242,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_254_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_254_inst_req_0;
      type_cast_254_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_254_inst_req_1;
      type_cast_254_inst_ack_1<= rack(0);
      type_cast_254_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_254_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call21_251,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv22_255,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_266_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_266_inst_req_0;
      type_cast_266_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_266_inst_req_1;
      type_cast_266_inst_ack_1<= rack(0);
      type_cast_266_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_266_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call25_263,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv28_267,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_279_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_279_inst_req_0;
      type_cast_279_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_279_inst_req_1;
      type_cast_279_inst_ack_1<= rack(0);
      type_cast_279_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_279_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call30_276,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv31_280,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_291_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_291_inst_req_0;
      type_cast_291_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_291_inst_req_1;
      type_cast_291_inst_ack_1<= rack(0);
      type_cast_291_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_291_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call34_288,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv37_292,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_304_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_304_inst_req_0;
      type_cast_304_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_304_inst_req_1;
      type_cast_304_inst_ack_1<= rack(0);
      type_cast_304_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_304_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call39_301,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv40_305,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_319_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_319_inst_req_0;
      type_cast_319_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_319_inst_req_1;
      type_cast_319_inst_ack_1<= rack(0);
      type_cast_319_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_319_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call44_316,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv47_320,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_332_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_332_inst_req_0;
      type_cast_332_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_332_inst_req_1;
      type_cast_332_inst_ack_1<= rack(0);
      type_cast_332_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_332_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call49_329,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv50_333,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_344_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_344_inst_req_0;
      type_cast_344_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_344_inst_req_1;
      type_cast_344_inst_ack_1<= rack(0);
      type_cast_344_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_344_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call53_341,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_345,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_357_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_357_inst_req_0;
      type_cast_357_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_357_inst_req_1;
      type_cast_357_inst_ack_1<= rack(0);
      type_cast_357_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_357_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call58_354,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv59_358,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_369_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_369_inst_req_0;
      type_cast_369_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_369_inst_req_1;
      type_cast_369_inst_ack_1<= rack(0);
      type_cast_369_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_369_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call62_366,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_370,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_382_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_382_inst_req_0;
      type_cast_382_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_382_inst_req_1;
      type_cast_382_inst_ack_1<= rack(0);
      type_cast_382_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_382_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call67_379,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv68_383,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_391_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_391_inst_req_0;
      type_cast_391_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_391_inst_req_1;
      type_cast_391_inst_ack_1<= rack(0);
      type_cast_391_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_391_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_260,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_392,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_395_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_395_inst_req_0;
      type_cast_395_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_395_inst_req_1;
      type_cast_395_inst_ack_1<= rack(0);
      type_cast_395_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_395_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add32_285,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_396,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_399_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_399_inst_req_0;
      type_cast_399_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_399_inst_req_1;
      type_cast_399_inst_ack_1<= rack(0);
      type_cast_399_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_399_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add41_310,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv77_400,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_420_inst
    process(sext_416) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := sext_416(63 downto 0);
      type_cast_420_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_425_inst
    process(ASHR_i64_i64_424_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_424_wire(63 downto 0);
      conv79_426 <= tmp_var; -- 
    end process;
    type_cast_467_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_467_inst_req_0;
      type_cast_467_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_467_inst_req_1;
      type_cast_467_inst_ack_1<= rack(0);
      type_cast_467_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_467_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_618,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_467_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_481_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_481_inst_req_0;
      type_cast_481_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_481_inst_req_1;
      type_cast_481_inst_ack_1<= rack(0);
      type_cast_481_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_481_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call85_478,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv86_482,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_494_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_494_inst_req_0;
      type_cast_494_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_494_inst_req_1;
      type_cast_494_inst_ack_1<= rack(0);
      type_cast_494_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_494_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call89_491,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv91_495,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_512_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_512_inst_req_0;
      type_cast_512_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_512_inst_req_1;
      type_cast_512_inst_ack_1<= rack(0);
      type_cast_512_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_512_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call95_509,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv97_513,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_530_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_530_inst_req_0;
      type_cast_530_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_530_inst_req_1;
      type_cast_530_inst_ack_1<= rack(0);
      type_cast_530_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_530_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call101_527,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv103_531,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_548_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_548_inst_req_0;
      type_cast_548_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_548_inst_req_1;
      type_cast_548_inst_ack_1<= rack(0);
      type_cast_548_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_548_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call107_545,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv109_549,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_566_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_566_inst_req_0;
      type_cast_566_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_566_inst_req_1;
      type_cast_566_inst_ack_1<= rack(0);
      type_cast_566_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_566_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call113_563,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv115_567,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_584_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_584_inst_req_0;
      type_cast_584_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_584_inst_req_1;
      type_cast_584_inst_ack_1<= rack(0);
      type_cast_584_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_584_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call119_581,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv121_585,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_602_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_602_inst_req_0;
      type_cast_602_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_602_inst_req_1;
      type_cast_602_inst_ack_1<= rack(0);
      type_cast_602_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_602_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call125_599,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv127_603,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_645_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_645_inst_req_0;
      type_cast_645_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_645_inst_req_1;
      type_cast_645_inst_ack_1<= rack(0);
      type_cast_645_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_645_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_644_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv179_646,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_649_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_649_inst_req_0;
      type_cast_649_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_649_inst_req_1;
      type_cast_649_inst_ack_1<= rack(0);
      type_cast_649_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_649_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add32_285,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv191_650,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_653_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_653_inst_req_0;
      type_cast_653_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_653_inst_req_1;
      type_cast_653_inst_ack_1<= rack(0);
      type_cast_653_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_653_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call43_313,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv193_654,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_668_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_668_inst_req_0;
      type_cast_668_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_668_inst_req_1;
      type_cast_668_inst_ack_1<= rack(0);
      type_cast_668_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_668_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_260,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv205_669,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_677_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_677_inst_req_0;
      type_cast_677_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_677_inst_req_1;
      type_cast_677_inst_ack_1<= rack(0);
      type_cast_677_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_677_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call43_313,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv240_678,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_712_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_712_inst_req_0;
      type_cast_712_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_712_inst_req_1;
      type_cast_712_inst_ack_1<= rack(0);
      type_cast_712_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_712_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => kx_x0_896,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_712_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_717_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_717_inst_req_0;
      type_cast_717_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_717_inst_req_1;
      type_cast_717_inst_ack_1<= rack(0);
      type_cast_717_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_717_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i138x_x1_924,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_717_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_722_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_722_inst_req_0;
      type_cast_722_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_722_inst_req_1;
      type_cast_722_inst_ack_1<= rack(0);
      type_cast_722_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_722_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x0_952,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_722_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_727_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_727_inst_req_0;
      type_cast_727_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_727_inst_req_1;
      type_cast_727_inst_ack_1<= rack(0);
      type_cast_727_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_727_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => kx_x1_709,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv177_728,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_731_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_731_inst_req_0;
      type_cast_731_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_731_inst_req_1;
      type_cast_731_inst_ack_1<= rack(0);
      type_cast_731_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_731_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv179_646,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_733_733_delayed_2_0_732,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_735_inst
    process(conv177_728) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv177_728(31 downto 0);
      type_cast_735_wire <= tmp_var; -- 
    end process;
    type_cast_778_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_778_inst_req_0;
      type_cast_778_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_778_inst_req_1;
      type_cast_778_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  ifx_xelse_exec_guard_764(0);
      type_cast_778_inst_gI: SplitGuardInterface generic map(name => "type_cast_778_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_778_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_778_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc187_774,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv189_779,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_795_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_795_inst_req_0;
      type_cast_795_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_795_inst_req_1;
      type_cast_795_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  ifx_xelse_exec_guard_777_delayed_1_0_791(0);
      type_cast_795_inst_gI: SplitGuardInterface generic map(name => "type_cast_795_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_795_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_795_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp196_788,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc201_796,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_829_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_829_inst_req_0;
      type_cast_829_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_829_inst_req_1;
      type_cast_829_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  ifx_xelse_exec_guard_796_delayed_2_0_825(0);
      type_cast_829_inst_gI: SplitGuardInterface generic map(name => "type_cast_829_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_829_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_829_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc201x_xi138x_x2_808,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv203_830,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_878_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_878_inst_req_0;
      type_cast_878_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_878_inst_req_1;
      type_cast_878_inst_ack_1<= rack(0);
      type_cast_878_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_878_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add184_758,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_834_834_delayed_3_0_879,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_902_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_902_inst_req_0;
      type_cast_902_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_902_inst_req_1;
      type_cast_902_inst_ack_1<= rack(0);
      type_cast_902_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_902_inst",
        buffer_size => 4,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i138x_x2_714,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_852_852_delayed_4_0_903,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_906_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_906_inst_req_0;
      type_cast_906_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_906_inst_req_1;
      type_cast_906_inst_ack_1<= rack(0);
      type_cast_906_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_906_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc201x_xi138x_x2_808,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_855_855_delayed_1_0_907,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_910_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_910_inst_req_0;
      type_cast_910_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_910_inst_req_1;
      type_cast_910_inst_ack_1<= rack(0);
      type_cast_910_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_910_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc201x_xi138x_x2_808,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_858_858_delayed_1_0_911,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_930_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_930_inst_req_0;
      type_cast_930_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_930_inst_req_1;
      type_cast_930_inst_ack_1<= rack(0);
      type_cast_930_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_930_inst",
        buffer_size => 4,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x1_719,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_868_868_delayed_4_0_931,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_934_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_934_inst_req_0;
      type_cast_934_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_934_inst_req_1;
      type_cast_934_inst_ack_1<= rack(0);
      type_cast_934_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_934_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x2_822,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_871_871_delayed_2_0_935,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_938_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_938_inst_req_0;
      type_cast_938_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_938_inst_req_1;
      type_cast_938_inst_ack_1<= rack(0);
      type_cast_938_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_938_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x2_822,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_874_874_delayed_2_0_939,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1212_index_1_rename
    process(R_idxprom290_1211_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom290_1211_resized;
      ov(13 downto 0) := iv;
      R_idxprom290_1211_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1212_index_1_resize
    process(idxprom290_1207) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom290_1207;
      ov := iv(13 downto 0);
      R_idxprom290_1211_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1212_root_address_inst
    process(array_obj_ref_1212_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1212_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1212_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1259_index_1_rename
    process(R_idxprom296_1258_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom296_1258_resized;
      ov(13 downto 0) := iv;
      R_idxprom296_1258_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1259_index_1_resize
    process(idxprom296_1254) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom296_1254;
      ov := iv(13 downto 0);
      R_idxprom296_1258_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1259_root_address_inst
    process(array_obj_ref_1259_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1259_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1259_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1305_index_1_rename
    process(R_idxprom302_1304_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom302_1304_resized;
      ov(13 downto 0) := iv;
      R_idxprom302_1304_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1305_index_1_resize
    process(idxprom302_1300) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom302_1300;
      ov := iv(13 downto 0);
      R_idxprom302_1304_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1305_root_address_inst
    process(array_obj_ref_1305_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1305_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1305_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_473_index_1_rename
    process(R_indvar_472_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_472_resized;
      ov(13 downto 0) := iv;
      R_indvar_472_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_473_index_1_resize
    process(indvar_461) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_461;
      ov := iv(13 downto 0);
      R_indvar_472_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_473_root_address_inst
    process(array_obj_ref_473_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_473_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_473_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1217_addr_0
    process(ptr_deref_1217_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1217_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1217_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1217_base_resize
    process(arrayidx291_1214) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx291_1214;
      ov := iv(13 downto 0);
      ptr_deref_1217_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1217_gather_scatter
    process(type_cast_1219_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_1219_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_1217_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1217_root_address_inst
    process(ptr_deref_1217_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1217_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1217_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1268_addr_0
    process(ptr_deref_1268_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1268_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1268_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1268_base_resize
    process(arrayidx297_1261) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx297_1261;
      ov := iv(13 downto 0);
      ptr_deref_1268_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1268_gather_scatter
    process(ptr_deref_1268_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1268_data_0;
      ov(63 downto 0) := iv;
      tmp298_1269 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1268_root_address_inst
    process(ptr_deref_1268_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1268_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1268_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1316_addr_0
    process(ptr_deref_1316_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1316_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1316_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1316_base_resize
    process(arrayidx303_1156_delayed_5_0_1313) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx303_1156_delayed_5_0_1313;
      ov := iv(13 downto 0);
      ptr_deref_1316_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1316_gather_scatter
    process(tmp298_1269) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp298_1269;
      ov(63 downto 0) := iv;
      ptr_deref_1316_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1316_root_address_inst
    process(ptr_deref_1316_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1316_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1316_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_610_addr_0
    process(ptr_deref_610_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_610_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_610_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_610_base_resize
    process(arrayidx_475) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_475;
      ov := iv(13 downto 0);
      ptr_deref_610_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_610_gather_scatter
    process(add128_608) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add128_608;
      ov(63 downto 0) := iv;
      ptr_deref_610_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_610_root_address_inst
    process(ptr_deref_610_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_610_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_610_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_707_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tobool_1324;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_707_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_707_branch_req_0,
          ack0 => do_while_stmt_707_branch_ack_0,
          ack1 => do_while_stmt_707_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1331_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ifx_xend304_whilex_xend_taken_1328;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1331_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1331_branch_req_0,
          ack0 => if_stmt_1331_branch_ack_0,
          ack1 => if_stmt_1331_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_433_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp390_432;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_433_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_433_branch_req_0,
          ack0 => if_stmt_433_branch_ack_0,
          ack1 => if_stmt_433_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_624_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond3_623;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_624_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_624_branch_req_0,
          ack0 => if_stmt_624_branch_ack_0,
          ack1 => if_stmt_624_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1021_inst
    process(sub241_1004, mul251_1016) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub241_1004, mul251_1016, tmp_var);
      tmp386_1022 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1033_inst
    process(tmp387_1028, kx_x0_896) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp387_1028, kx_x0_896, tmp_var);
      add252_1034 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_640_inst
    process(add41_310) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add41_310, type_cast_639_wire_constant, tmp_var);
      sub_641 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_757_inst
    process(kx_x1_748_delayed_1_0_751) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(kx_x1_748_delayed_1_0_751, type_cast_756_wire_constant, tmp_var);
      add184_758 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_773_inst
    process(jx_x1_761_delayed_1_0_767) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(jx_x1_761_delayed_1_0_767, type_cast_772_wire_constant, tmp_var);
      inc187_774 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_807_inst
    process(inc201_796, i138x_x2_785_delayed_3_0_802) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc201_796, i138x_x2_785_delayed_3_0_802, tmp_var);
      inc201x_xi138x_x2_808 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_985_inst
    process(jx_x0_952, mul229_980) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(jx_x0_952, mul229_980, tmp_var);
      tmp_986 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_997_inst
    process(tmp385_992, kx_x0_896) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp385_992, kx_x0_896, tmp_var);
      add230_998 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_664_inst
    process(shl194_660, conv191_650) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl194_660, conv191_650, tmp_var);
      add195_665 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_673_inst
    process(shl194_660, conv205_669) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl194_660, conv205_669, tmp_var);
      add209_674 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_682_inst
    process(conv193_654, conv205_669) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv193_654, conv205_669, tmp_var);
      add266_683 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_687_inst
    process(conv193_654, conv191_650) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv193_654, conv191_650, tmp_var);
      add283_688 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_617_inst
    process(indvar_461) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_461, type_cast_616_wire_constant, tmp_var);
      indvarx_xnext_618 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1080_inst
    process(cmp258x_xnot_1058, cmp267_1072) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmp258x_xnot_1058, cmp267_1072, tmp_var);
      orx_xcond_1081 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1088_inst
    process(ifx_xend214_exec_guard_993_delayed_1_0_1084, orx_xcond_1081) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(ifx_xend214_exec_guard_993_delayed_1_0_1084, orx_xcond_1081, tmp_var);
      ifx_xend214_lorx_xlhsx_xfalse269_taken_1089 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1097_inst
    process(ifx_xend214_exec_guard_998_delayed_1_0_1092, NOT_u1_u1_1096_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(ifx_xend214_exec_guard_998_delayed_1_0_1092, NOT_u1_u1_1096_wire, tmp_var);
      ifx_xend214_ifx_xthen286_taken_1098 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1150_inst
    process(cmp274x_xnot_1128, cmp284_1142) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmp274x_xnot_1128, cmp284_1142, tmp_var);
      orx_xcond393_1151 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1158_inst
    process(lorx_xlhsx_xfalse269_exec_guard_1039_delayed_1_0_1154, orx_xcond393_1151) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(lorx_xlhsx_xfalse269_exec_guard_1039_delayed_1_0_1154, orx_xcond393_1151, tmp_var);
      lorx_xlhsx_xfalse269_ifx_xelse292_taken_1159 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1167_inst
    process(lorx_xlhsx_xfalse269_exec_guard_1044_delayed_1_0_1162, NOT_u1_u1_1166_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(lorx_xlhsx_xfalse269_exec_guard_1044_delayed_1_0_1162, NOT_u1_u1_1166_wire, tmp_var);
      lorx_xlhsx_xfalse269_ifx_xthen286_taken_1168 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_846_inst
    process(ifx_xelse_exec_guard_808_delayed_3_0_842, cmp210_839) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(ifx_xelse_exec_guard_808_delayed_3_0_842, cmp210_839, tmp_var);
      ifx_xelse_ifx_xthen212_taken_847 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_855_inst
    process(ifx_xelse_exec_guard_813_delayed_3_0_850, NOT_u1_u1_854_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(ifx_xelse_exec_guard_813_delayed_3_0_850, NOT_u1_u1_854_wire, tmp_var);
      ifx_xelse_ifx_xend214_taken_856 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1196_inst
    process(type_cast_1192_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1192_wire, type_cast_1195_wire_constant, tmp_var);
      ASHR_i32_i32_1196_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1243_inst
    process(type_cast_1239_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1239_wire, type_cast_1242_wire_constant, tmp_var);
      ASHR_i32_i32_1243_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1289_inst
    process(type_cast_1285_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1285_wire, type_cast_1288_wire_constant, tmp_var);
      ASHR_i32_i32_1289_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_424_inst
    process(type_cast_420_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_420_wire, type_cast_423_wire_constant, tmp_var);
      ASHR_i64_i64_424_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1323_inst
    process(flagx_x0_974) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(flagx_x0_974, type_cast_1322_wire_constant, tmp_var);
      tobool_1324 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_787_inst
    process(conv189_779, add195_665) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv189_779, add195_665, tmp_var);
      cmp196_788 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_838_inst
    process(conv203_830, add209_674) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv203_830, add209_674, tmp_var);
      cmp210_839 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_622_inst
    process(indvarx_xnext_618, umax2_458) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_618, umax2_458, tmp_var);
      exitcond3_623 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1362_inst
    process(sub314_1353) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub314_1353, type_cast_1361_wire_constant, tmp_var);
      shr320_1363 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1372_inst
    process(sub314_1353) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub314_1353, type_cast_1371_wire_constant, tmp_var);
      shr326_1373 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1382_inst
    process(sub314_1353) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub314_1353, type_cast_1381_wire_constant, tmp_var);
      shr332_1383 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1392_inst
    process(sub314_1353) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub314_1353, type_cast_1391_wire_constant, tmp_var);
      shr338_1393 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1402_inst
    process(sub314_1353) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub314_1353, type_cast_1401_wire_constant, tmp_var);
      shr344_1403 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1412_inst
    process(sub314_1353) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub314_1353, type_cast_1411_wire_constant, tmp_var);
      shr350_1413 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1422_inst
    process(sub314_1353) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub314_1353, type_cast_1421_wire_constant, tmp_var);
      shr356_1423 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_444_inst
    process(conv79_426) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv79_426, type_cast_443_wire_constant, tmp_var);
      shr_445 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1015_inst
    process(add32_285, sub250_1010) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(add32_285, sub250_1010, tmp_var);
      mul251_1016 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1027_inst
    process(tmp386_1022, add41_310) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp386_1022, add41_310, tmp_var);
      tmp387_1028 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_979_inst
    process(add60_363, i138x_x1_924) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(add60_363, i138x_x1_924, tmp_var);
      mul229_980 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_991_inst
    process(tmp_986, add69_388) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp_986, add69_388, tmp_var);
      tmp385_992 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1464_inst
    process(conv380_1456, add51_338) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv380_1456, add51_338, tmp_var);
      mul381_1465 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1469_inst
    process(mul381_1465, conv383_1460) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul381_1465, conv383_1460, tmp_var);
      mul384_1470 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_410_inst
    process(mul_406, conv75_396) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_406, conv75_396, tmp_var);
      mul78_411 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_415_inst
    process(mul78_411, conv77_400) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul78_411, conv77_400, tmp_var);
      sext_416 <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1096_inst
    process(orx_xcond_1081) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", orx_xcond_1081, tmp_var);
      NOT_u1_u1_1096_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1166_inst
    process(orx_xcond393_1151) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", orx_xcond393_1151, tmp_var);
      NOT_u1_u1_1166_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1327_inst
    process(tobool_1324) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", tobool_1324, tmp_var);
      ifx_xend304_whilex_xend_taken_1328 <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_744_inst
    process(cmp180_738) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp180_738, tmp_var);
      whilex_xbody_ifx_xthen_taken_745 <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_854_inst
    process(cmp210_839) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp210_839, tmp_var);
      NOT_u1_u1_854_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u16_u16_259_inst
    process(shl20_248, conv22_255) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl20_248, conv22_255, tmp_var);
      add23_260 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_284_inst
    process(shl29_273, conv31_280) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl29_273, conv31_280, tmp_var);
      add32_285 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_309_inst
    process(shl38_298, conv40_305) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl38_298, conv40_305, tmp_var);
      add41_310 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_362_inst
    process(shl57_351, conv59_358) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl57_351, conv59_358, tmp_var);
      add60_363 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_387_inst
    process(shl66_376, conv68_383) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl66_376, conv68_383, tmp_var);
      add69_388 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1175_inst
    process(ifx_xend214_ifx_xthen286_taken_1050_delayed_1_0_1171, lorx_xlhsx_xfalse269_ifx_xthen286_taken_1168) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(ifx_xend214_ifx_xthen286_taken_1050_delayed_1_0_1171, lorx_xlhsx_xfalse269_ifx_xthen286_taken_1168, tmp_var);
      ifx_xthen286_exec_guard_1176 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_870_inst
    process(ifx_xthen_ifx_xend214_taken_826_delayed_3_0_865, ifx_xthen212_ifx_xend214_taken_862) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(ifx_xthen_ifx_xend214_taken_826_delayed_3_0_865, ifx_xthen212_ifx_xend214_taken_862, tmp_var);
      OR_u1_u1_870_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_871_inst
    process(ifx_xelse_ifx_xend214_taken_856, OR_u1_u1_870_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(ifx_xelse_ifx_xend214_taken_856, OR_u1_u1_870_wire, tmp_var);
      ifx_xend214_exec_guard_872 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_337_inst
    process(shl48_326, conv50_333) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl48_326, conv50_333, tmp_var);
      add51_338 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_499_inst
    process(shl88_488, conv91_495) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl88_488, conv91_495, tmp_var);
      add92_500 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_517_inst
    process(shl94_506, conv97_513) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl94_506, conv97_513, tmp_var);
      add98_518 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_535_inst
    process(shl100_524, conv103_531) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl100_524, conv103_531, tmp_var);
      add104_536 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_553_inst
    process(shl106_542, conv109_549) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl106_542, conv109_549, tmp_var);
      add110_554 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_571_inst
    process(shl112_560, conv115_567) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl112_560, conv115_567, tmp_var);
      add116_572 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_589_inst
    process(shl118_578, conv121_585) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl118_578, conv121_585, tmp_var);
      add122_590 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_607_inst
    process(shl124_596, conv127_603) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl124_596, conv127_603, tmp_var);
      add128_608 <= tmp_var; --
    end process;
    -- binary operator SGT_i32_u1_737_inst
    process(type_cast_735_wire, type_cast_733_733_delayed_2_0_732) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(type_cast_735_wire, type_cast_733_733_delayed_2_0_732, tmp_var);
      cmp180_738 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_247_inst
    process(conv19_242) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv19_242, type_cast_246_wire_constant, tmp_var);
      shl20_248 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_272_inst
    process(conv28_267) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv28_267, type_cast_271_wire_constant, tmp_var);
      shl29_273 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_297_inst
    process(conv37_292) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv37_292, type_cast_296_wire_constant, tmp_var);
      shl38_298 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_350_inst
    process(conv56_345) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv56_345, type_cast_349_wire_constant, tmp_var);
      shl57_351 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_375_inst
    process(conv65_370) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv65_370, type_cast_374_wire_constant, tmp_var);
      shl66_376 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_325_inst
    process(conv47_320) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv47_320, type_cast_324_wire_constant, tmp_var);
      shl48_326 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_659_inst
    process(conv193_654) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv193_654, type_cast_658_wire_constant, tmp_var);
      shl194_660 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_405_inst
    process(conv73_392) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv73_392, type_cast_404_wire_constant, tmp_var);
      mul_406 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_487_inst
    process(conv86_482) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv86_482, type_cast_486_wire_constant, tmp_var);
      shl88_488 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_505_inst
    process(add92_500) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add92_500, type_cast_504_wire_constant, tmp_var);
      shl94_506 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_523_inst
    process(add98_518) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add98_518, type_cast_522_wire_constant, tmp_var);
      shl100_524 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_541_inst
    process(add104_536) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add104_536, type_cast_540_wire_constant, tmp_var);
      shl106_542 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_559_inst
    process(add110_554) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add110_554, type_cast_558_wire_constant, tmp_var);
      shl112_560 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_577_inst
    process(add116_572) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add116_572, type_cast_576_wire_constant, tmp_var);
      shl118_578 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_595_inst
    process(add122_590) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add122_590, type_cast_594_wire_constant, tmp_var);
      shl124_596 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1071_inst
    process(type_cast_1069_wire, type_cast_983_983_delayed_1_0_1065) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1069_wire, type_cast_983_983_delayed_1_0_1065, tmp_var);
      cmp267_1072 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1141_inst
    process(type_cast_1139_wire, type_cast_1029_1029_delayed_1_0_1135) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1139_wire, type_cast_1029_1029_delayed_1_0_1135, tmp_var);
      cmp284_1142 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1003_inst
    process(jx_x0_952, conv240_678) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(jx_x0_952, conv240_678, tmp_var);
      sub241_1004 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1009_inst
    process(i138x_x1_924, conv240_678) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(i138x_x1_924, conv240_678, tmp_var);
      sub250_1010 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_1352_inst
    process(conv310_1348, conv134_1340) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv310_1348, conv134_1340, tmp_var);
      sub314_1353 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_431_inst
    process(conv79_426) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(conv79_426, type_cast_430_wire_constant, tmp_var);
      cmp390_432 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_450_inst
    process(shr_445) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(shr_445, type_cast_449_wire_constant, tmp_var);
      tmp1_451 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1047_inst
    process(conv255_1039, conv193_654) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(conv255_1039, conv193_654, tmp_var);
      cmp258_1048 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1117_inst
    process(conv271_1109, conv193_654) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(conv271_1109, conv193_654, tmp_var);
      cmp274_1118 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_1057_inst
    process(cmp258_1048) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp258_1048, type_cast_1056_wire_constant, tmp_var);
      cmp258x_xnot_1058 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_1127_inst
    process(cmp274_1118) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp274_1118, type_cast_1126_wire_constant, tmp_var);
      cmp274x_xnot_1128 <= tmp_var; --
    end process;
    -- shared split operator group (93) : array_obj_ref_1212_index_offset 
    ApIntAdd_group_93: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom290_1211_scaled;
      array_obj_ref_1212_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1212_index_offset_req_0;
      array_obj_ref_1212_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1212_index_offset_req_1;
      array_obj_ref_1212_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_93_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_93_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_93",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 93
    -- shared split operator group (94) : array_obj_ref_1259_index_offset 
    ApIntAdd_group_94: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom296_1258_scaled;
      array_obj_ref_1259_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1259_index_offset_req_0;
      array_obj_ref_1259_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1259_index_offset_req_1;
      array_obj_ref_1259_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_94_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_94_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_94",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 94
    -- shared split operator group (95) : array_obj_ref_1305_index_offset 
    ApIntAdd_group_95: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom302_1304_scaled;
      array_obj_ref_1305_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1305_index_offset_req_0;
      array_obj_ref_1305_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1305_index_offset_req_1;
      array_obj_ref_1305_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_95_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_95_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_95",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 95
    -- shared split operator group (96) : array_obj_ref_473_index_offset 
    ApIntAdd_group_96: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_472_scaled;
      array_obj_ref_473_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_473_index_offset_req_0;
      array_obj_ref_473_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_473_index_offset_req_1;
      array_obj_ref_473_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_96_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_96_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_96",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 96
    -- unary operator type_cast_1183_inst
    process(add230_1056_delayed_2_0_1179) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", add230_1056_delayed_2_0_1179, tmp_var);
      type_cast_1183_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1205_inst
    process(shr289_1198) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr289_1198, tmp_var);
      type_cast_1205_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1230_inst
    process(add252_1094_delayed_2_0_1226) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", add252_1094_delayed_2_0_1226, tmp_var);
      type_cast_1230_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1252_inst
    process(shr295_1245) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr295_1245, tmp_var);
      type_cast_1252_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1276_inst
    process(add230_1128_delayed_2_0_1272) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", add230_1128_delayed_2_0_1272, tmp_var);
      type_cast_1276_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1298_inst
    process(shr301_1291) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr301_1291, tmp_var);
      type_cast_1298_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1338_inst
    process(call133_635) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call133_635, tmp_var);
      type_cast_1338_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1346_inst
    process(call309_1343) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call309_1343, tmp_var);
      type_cast_1346_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_644_inst
    process(sub_641) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", sub_641, tmp_var);
      type_cast_644_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_1268_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1268_load_0_req_0;
      ptr_deref_1268_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1268_load_0_req_1;
      ptr_deref_1268_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= ifx_xelse292_exec_guard_1121_delayed_8_0_1264(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1268_word_address_0;
      ptr_deref_1268_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_1316_store_0 ptr_deref_1217_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 2, 0 => 2);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 15, 0 => 15);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => true, 1 => true);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 6, 1 => 6);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1316_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1217_store_0_req_0;
      ptr_deref_1316_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1217_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1316_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1217_store_0_req_1;
      ptr_deref_1316_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1217_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= ifx_xthen286_exec_guard_1176(0);
      guard_vector(1)  <= ifx_xelse292_exec_guard_1155_delayed_14_0_1310(0);
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1316_word_address_0 & ptr_deref_1217_word_address_0;
      data_in <= ptr_deref_1316_data_0 & ptr_deref_1217_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_610_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_610_store_0_req_0;
      ptr_deref_610_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_610_store_0_req_1;
      ptr_deref_610_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_610_word_address_0;
      data_in <= ptr_deref_610_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared inport operator group (0) : RPIPE_zeropad_input_pipe_275_inst RPIPE_zeropad_input_pipe_236_inst RPIPE_zeropad_input_pipe_233_inst RPIPE_zeropad_input_pipe_230_inst RPIPE_zeropad_input_pipe_262_inst RPIPE_zeropad_input_pipe_227_inst RPIPE_zeropad_input_pipe_224_inst RPIPE_zeropad_input_pipe_287_inst RPIPE_zeropad_input_pipe_250_inst RPIPE_zeropad_input_pipe_328_inst RPIPE_zeropad_input_pipe_378_inst RPIPE_zeropad_input_pipe_365_inst RPIPE_zeropad_input_pipe_300_inst RPIPE_zeropad_input_pipe_315_inst RPIPE_zeropad_input_pipe_340_inst RPIPE_zeropad_input_pipe_353_inst RPIPE_zeropad_input_pipe_312_inst RPIPE_zeropad_input_pipe_477_inst RPIPE_zeropad_input_pipe_490_inst RPIPE_zeropad_input_pipe_508_inst RPIPE_zeropad_input_pipe_526_inst RPIPE_zeropad_input_pipe_544_inst RPIPE_zeropad_input_pipe_562_inst RPIPE_zeropad_input_pipe_580_inst RPIPE_zeropad_input_pipe_598_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(199 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 24 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 24 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 24 downto 0);
      signal guard_vector : std_logic_vector( 24 downto 0);
      constant outBUFs : IntegerArray(24 downto 0) := (24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(24 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false);
      constant guardBuffering: IntegerArray(24 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2);
      -- 
    begin -- 
      reqL_unguarded(24) <= RPIPE_zeropad_input_pipe_275_inst_req_0;
      reqL_unguarded(23) <= RPIPE_zeropad_input_pipe_236_inst_req_0;
      reqL_unguarded(22) <= RPIPE_zeropad_input_pipe_233_inst_req_0;
      reqL_unguarded(21) <= RPIPE_zeropad_input_pipe_230_inst_req_0;
      reqL_unguarded(20) <= RPIPE_zeropad_input_pipe_262_inst_req_0;
      reqL_unguarded(19) <= RPIPE_zeropad_input_pipe_227_inst_req_0;
      reqL_unguarded(18) <= RPIPE_zeropad_input_pipe_224_inst_req_0;
      reqL_unguarded(17) <= RPIPE_zeropad_input_pipe_287_inst_req_0;
      reqL_unguarded(16) <= RPIPE_zeropad_input_pipe_250_inst_req_0;
      reqL_unguarded(15) <= RPIPE_zeropad_input_pipe_328_inst_req_0;
      reqL_unguarded(14) <= RPIPE_zeropad_input_pipe_378_inst_req_0;
      reqL_unguarded(13) <= RPIPE_zeropad_input_pipe_365_inst_req_0;
      reqL_unguarded(12) <= RPIPE_zeropad_input_pipe_300_inst_req_0;
      reqL_unguarded(11) <= RPIPE_zeropad_input_pipe_315_inst_req_0;
      reqL_unguarded(10) <= RPIPE_zeropad_input_pipe_340_inst_req_0;
      reqL_unguarded(9) <= RPIPE_zeropad_input_pipe_353_inst_req_0;
      reqL_unguarded(8) <= RPIPE_zeropad_input_pipe_312_inst_req_0;
      reqL_unguarded(7) <= RPIPE_zeropad_input_pipe_477_inst_req_0;
      reqL_unguarded(6) <= RPIPE_zeropad_input_pipe_490_inst_req_0;
      reqL_unguarded(5) <= RPIPE_zeropad_input_pipe_508_inst_req_0;
      reqL_unguarded(4) <= RPIPE_zeropad_input_pipe_526_inst_req_0;
      reqL_unguarded(3) <= RPIPE_zeropad_input_pipe_544_inst_req_0;
      reqL_unguarded(2) <= RPIPE_zeropad_input_pipe_562_inst_req_0;
      reqL_unguarded(1) <= RPIPE_zeropad_input_pipe_580_inst_req_0;
      reqL_unguarded(0) <= RPIPE_zeropad_input_pipe_598_inst_req_0;
      RPIPE_zeropad_input_pipe_275_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_zeropad_input_pipe_236_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_zeropad_input_pipe_233_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_zeropad_input_pipe_230_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_zeropad_input_pipe_262_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_zeropad_input_pipe_227_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_zeropad_input_pipe_224_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_zeropad_input_pipe_287_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_zeropad_input_pipe_250_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_zeropad_input_pipe_328_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_zeropad_input_pipe_378_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_zeropad_input_pipe_365_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_zeropad_input_pipe_300_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_zeropad_input_pipe_315_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_zeropad_input_pipe_340_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_zeropad_input_pipe_353_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_zeropad_input_pipe_312_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_zeropad_input_pipe_477_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_zeropad_input_pipe_490_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_zeropad_input_pipe_508_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_zeropad_input_pipe_526_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_zeropad_input_pipe_544_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_zeropad_input_pipe_562_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_zeropad_input_pipe_580_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_zeropad_input_pipe_598_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(24) <= RPIPE_zeropad_input_pipe_275_inst_req_1;
      reqR_unguarded(23) <= RPIPE_zeropad_input_pipe_236_inst_req_1;
      reqR_unguarded(22) <= RPIPE_zeropad_input_pipe_233_inst_req_1;
      reqR_unguarded(21) <= RPIPE_zeropad_input_pipe_230_inst_req_1;
      reqR_unguarded(20) <= RPIPE_zeropad_input_pipe_262_inst_req_1;
      reqR_unguarded(19) <= RPIPE_zeropad_input_pipe_227_inst_req_1;
      reqR_unguarded(18) <= RPIPE_zeropad_input_pipe_224_inst_req_1;
      reqR_unguarded(17) <= RPIPE_zeropad_input_pipe_287_inst_req_1;
      reqR_unguarded(16) <= RPIPE_zeropad_input_pipe_250_inst_req_1;
      reqR_unguarded(15) <= RPIPE_zeropad_input_pipe_328_inst_req_1;
      reqR_unguarded(14) <= RPIPE_zeropad_input_pipe_378_inst_req_1;
      reqR_unguarded(13) <= RPIPE_zeropad_input_pipe_365_inst_req_1;
      reqR_unguarded(12) <= RPIPE_zeropad_input_pipe_300_inst_req_1;
      reqR_unguarded(11) <= RPIPE_zeropad_input_pipe_315_inst_req_1;
      reqR_unguarded(10) <= RPIPE_zeropad_input_pipe_340_inst_req_1;
      reqR_unguarded(9) <= RPIPE_zeropad_input_pipe_353_inst_req_1;
      reqR_unguarded(8) <= RPIPE_zeropad_input_pipe_312_inst_req_1;
      reqR_unguarded(7) <= RPIPE_zeropad_input_pipe_477_inst_req_1;
      reqR_unguarded(6) <= RPIPE_zeropad_input_pipe_490_inst_req_1;
      reqR_unguarded(5) <= RPIPE_zeropad_input_pipe_508_inst_req_1;
      reqR_unguarded(4) <= RPIPE_zeropad_input_pipe_526_inst_req_1;
      reqR_unguarded(3) <= RPIPE_zeropad_input_pipe_544_inst_req_1;
      reqR_unguarded(2) <= RPIPE_zeropad_input_pipe_562_inst_req_1;
      reqR_unguarded(1) <= RPIPE_zeropad_input_pipe_580_inst_req_1;
      reqR_unguarded(0) <= RPIPE_zeropad_input_pipe_598_inst_req_1;
      RPIPE_zeropad_input_pipe_275_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_zeropad_input_pipe_236_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_zeropad_input_pipe_233_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_zeropad_input_pipe_230_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_zeropad_input_pipe_262_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_zeropad_input_pipe_227_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_zeropad_input_pipe_224_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_zeropad_input_pipe_287_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_zeropad_input_pipe_250_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_zeropad_input_pipe_328_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_zeropad_input_pipe_378_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_zeropad_input_pipe_365_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_zeropad_input_pipe_300_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_zeropad_input_pipe_315_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_zeropad_input_pipe_340_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_zeropad_input_pipe_353_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_zeropad_input_pipe_312_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_zeropad_input_pipe_477_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_zeropad_input_pipe_490_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_zeropad_input_pipe_508_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_zeropad_input_pipe_526_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_zeropad_input_pipe_544_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_zeropad_input_pipe_562_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_zeropad_input_pipe_580_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_zeropad_input_pipe_598_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      call30_276 <= data_out(199 downto 192);
      call16_237 <= data_out(191 downto 184);
      call11_234 <= data_out(183 downto 176);
      call6_231 <= data_out(175 downto 168);
      call25_263 <= data_out(167 downto 160);
      call2_228 <= data_out(159 downto 152);
      call_225 <= data_out(151 downto 144);
      call34_288 <= data_out(143 downto 136);
      call21_251 <= data_out(135 downto 128);
      call49_329 <= data_out(127 downto 120);
      call67_379 <= data_out(119 downto 112);
      call62_366 <= data_out(111 downto 104);
      call39_301 <= data_out(103 downto 96);
      call44_316 <= data_out(95 downto 88);
      call53_341 <= data_out(87 downto 80);
      call58_354 <= data_out(79 downto 72);
      call43_313 <= data_out(71 downto 64);
      call85_478 <= data_out(63 downto 56);
      call89_491 <= data_out(55 downto 48);
      call95_509 <= data_out(47 downto 40);
      call101_527 <= data_out(39 downto 32);
      call107_545 <= data_out(31 downto 24);
      call113_563 <= data_out(23 downto 16);
      call119_581 <= data_out(15 downto 8);
      call125_599 <= data_out(7 downto 0);
      zeropad_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "zeropad_input_pipe_read_0_gI", nreqs => 25, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      zeropad_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "zeropad_input_pipe_read_0", data_width => 8,  num_reqs => 25,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => zeropad_input_pipe_pipe_read_req(0),
          oack => zeropad_input_pipe_pipe_read_ack(0),
          odata => zeropad_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_zeropad_output_pipe_1434_inst WPIPE_zeropad_output_pipe_1446_inst WPIPE_zeropad_output_pipe_1440_inst WPIPE_zeropad_output_pipe_1431_inst WPIPE_zeropad_output_pipe_1443_inst WPIPE_zeropad_output_pipe_1437_inst WPIPE_zeropad_output_pipe_1428_inst WPIPE_zeropad_output_pipe_1449_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 7 downto 0);
      signal update_req, update_ack : BooleanArray( 7 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 7 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      sample_req_unguarded(7) <= WPIPE_zeropad_output_pipe_1434_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_zeropad_output_pipe_1446_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_zeropad_output_pipe_1440_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_zeropad_output_pipe_1431_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_zeropad_output_pipe_1443_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_zeropad_output_pipe_1437_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_zeropad_output_pipe_1428_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_zeropad_output_pipe_1449_inst_req_0;
      WPIPE_zeropad_output_pipe_1434_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_zeropad_output_pipe_1446_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_zeropad_output_pipe_1440_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_zeropad_output_pipe_1431_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_zeropad_output_pipe_1443_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_zeropad_output_pipe_1437_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_zeropad_output_pipe_1428_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_zeropad_output_pipe_1449_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(7) <= WPIPE_zeropad_output_pipe_1434_inst_req_1;
      update_req_unguarded(6) <= WPIPE_zeropad_output_pipe_1446_inst_req_1;
      update_req_unguarded(5) <= WPIPE_zeropad_output_pipe_1440_inst_req_1;
      update_req_unguarded(4) <= WPIPE_zeropad_output_pipe_1431_inst_req_1;
      update_req_unguarded(3) <= WPIPE_zeropad_output_pipe_1443_inst_req_1;
      update_req_unguarded(2) <= WPIPE_zeropad_output_pipe_1437_inst_req_1;
      update_req_unguarded(1) <= WPIPE_zeropad_output_pipe_1428_inst_req_1;
      update_req_unguarded(0) <= WPIPE_zeropad_output_pipe_1449_inst_req_1;
      WPIPE_zeropad_output_pipe_1434_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_zeropad_output_pipe_1446_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_zeropad_output_pipe_1440_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_zeropad_output_pipe_1431_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_zeropad_output_pipe_1443_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_zeropad_output_pipe_1437_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_zeropad_output_pipe_1428_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_zeropad_output_pipe_1449_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      data_in <= conv347_1407 & conv323_1367 & conv335_1387 & conv353_1417 & conv329_1377 & conv341_1397 & conv359_1427 & conv317_1357;
      zeropad_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "zeropad_output_pipe_write_0_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      zeropad_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "zeropad_output_pipe", data_width => 8, num_reqs => 8, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => zeropad_output_pipe_pipe_write_req(0),
          oack => zeropad_output_pipe_pipe_write_ack(0),
          odata => zeropad_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_1343_call call_stmt_635_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_1343_call_req_0;
      reqL_unguarded(0) <= call_stmt_635_call_req_0;
      call_stmt_1343_call_ack_0 <= ackL_unguarded(1);
      call_stmt_635_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_1343_call_req_1;
      reqR_unguarded(0) <= call_stmt_635_call_req_1;
      call_stmt_1343_call_ack_1 <= ackR_unguarded(1);
      call_stmt_635_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call309_1343 <= data_out(127 downto 64);
      call133_635 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1472_call 
    sendOutput_call_group_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1472_call_req_0;
      call_stmt_1472_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1472_call_req_1;
      call_stmt_1472_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      sendOutput_call_group_1_gI: SplitGuardInterface generic map(name => "sendOutput_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= mul384_1470;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 32,
        owidth => 32,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => sendOutput_call_reqs(0),
          ackR => sendOutput_call_acks(0),
          dataR => sendOutput_call_data(31 downto 0),
          tagR => sendOutput_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => sendOutput_return_acks(0), -- cross-over
          ackL => sendOutput_return_reqs(0), -- cross-over
          tagL => sendOutput_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end zeropad3D_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    zeropad_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    zeropad_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    zeropad_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    zeropad_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(17 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(17 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(0 downto 0);
  -- declarations related to module sendOutput
  component sendOutput is -- 
    generic (tag_length : integer); 
    port ( -- 
      size : in  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      zeropad_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module sendOutput
  signal sendOutput_size :  std_logic_vector(31 downto 0);
  signal sendOutput_in_args    : std_logic_vector(31 downto 0);
  signal sendOutput_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal sendOutput_tag_out   : std_logic_vector(1 downto 0);
  signal sendOutput_start_req : std_logic;
  signal sendOutput_start_ack : std_logic;
  signal sendOutput_fin_req   : std_logic;
  signal sendOutput_fin_ack : std_logic;
  -- caller side aggregated signals for module sendOutput
  signal sendOutput_call_reqs: std_logic_vector(0 downto 0);
  signal sendOutput_call_acks: std_logic_vector(0 downto 0);
  signal sendOutput_return_reqs: std_logic_vector(0 downto 0);
  signal sendOutput_return_acks: std_logic_vector(0 downto 0);
  signal sendOutput_call_data: std_logic_vector(31 downto 0);
  signal sendOutput_call_tag: std_logic_vector(0 downto 0);
  signal sendOutput_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_c :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module timerDaemon
  component timerDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timerDaemon
  signal timerDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal timerDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal timerDaemon_start_req : std_logic;
  signal timerDaemon_start_ack : std_logic;
  signal timerDaemon_fin_req   : std_logic;
  signal timerDaemon_fin_ack : std_logic;
  -- declarations related to module zeropad3D
  component zeropad3D is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      zeropad_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      zeropad_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      zeropad_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      zeropad_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      sendOutput_call_reqs : out  std_logic_vector(0 downto 0);
      sendOutput_call_acks : in   std_logic_vector(0 downto 0);
      sendOutput_call_data : out  std_logic_vector(31 downto 0);
      sendOutput_call_tag  :  out  std_logic_vector(0 downto 0);
      sendOutput_return_reqs : out  std_logic_vector(0 downto 0);
      sendOutput_return_acks : in   std_logic_vector(0 downto 0);
      sendOutput_return_tag :  in   std_logic_vector(0 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module zeropad3D
  signal zeropad3D_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal zeropad3D_tag_out   : std_logic_vector(1 downto 0);
  signal zeropad3D_start_req : std_logic;
  signal zeropad3D_start_ack : std_logic;
  signal zeropad3D_fin_req   : std_logic;
  signal zeropad3D_fin_ack : std_logic;
  -- aggregate signals for read from pipe zeropad_input_pipe
  signal zeropad_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal zeropad_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal zeropad_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe zeropad_output_pipe
  signal zeropad_output_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal zeropad_output_pipe_pipe_write_req: std_logic_vector(1 downto 0);
  signal zeropad_output_pipe_pipe_write_ack: std_logic_vector(1 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module sendOutput
  sendOutput_size <= sendOutput_in_args(31 downto 0);
  -- call arbiter for module sendOutput
  sendOutput_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 32,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => sendOutput_call_reqs,
      call_acks => sendOutput_call_acks,
      return_reqs => sendOutput_return_reqs,
      return_acks => sendOutput_return_acks,
      call_data  => sendOutput_call_data,
      call_tag  => sendOutput_call_tag,
      return_tag  => sendOutput_return_tag,
      call_mtag => sendOutput_tag_in,
      return_mtag => sendOutput_tag_out,
      call_mreq => sendOutput_start_req,
      call_mack => sendOutput_start_ack,
      return_mreq => sendOutput_fin_req,
      return_mack => sendOutput_fin_ack,
      call_mdata => sendOutput_in_args,
      clk => clk, 
      reset => reset --
    ); --
  sendOutput_instance:sendOutput-- 
    generic map(tag_length => 2)
    port map(-- 
      size => sendOutput_size,
      start_req => sendOutput_start_req,
      start_ack => sendOutput_start_ack,
      fin_req => sendOutput_fin_req,
      fin_ack => sendOutput_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(18 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(1 downto 0),
      zeropad_output_pipe_pipe_write_req => zeropad_output_pipe_pipe_write_req(1 downto 1),
      zeropad_output_pipe_pipe_write_ack => zeropad_output_pipe_pipe_write_ack(1 downto 1),
      zeropad_output_pipe_pipe_write_data => zeropad_output_pipe_pipe_write_data(15 downto 8),
      tag_in => sendOutput_tag_in,
      tag_out => sendOutput_tag_out-- 
    ); -- 
  -- module timer
  timer_out_args <= timer_c ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      c => timer_c,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(0 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(17 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  -- module timerDaemon
  timerDaemon_instance:timerDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => timerDaemon_start_req,
      start_ack => timerDaemon_start_ack,
      fin_req => timerDaemon_fin_req,
      fin_ack => timerDaemon_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(0 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(63 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(17 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(0 downto 0),
      tag_in => timerDaemon_tag_in,
      tag_out => timerDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  timerDaemon_tag_in <= (others => '0');
  timerDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => timerDaemon_start_req, start_ack => timerDaemon_start_ack,  fin_req => timerDaemon_fin_req,  fin_ack => timerDaemon_fin_ack);
  -- module zeropad3D
  zeropad3D_instance:zeropad3D-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => zeropad3D_start_req,
      start_ack => zeropad3D_start_ack,
      fin_req => zeropad3D_fin_req,
      fin_ack => zeropad3D_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(17 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(0 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(13 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(18 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(1 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(17 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(0 downto 0),
      zeropad_input_pipe_pipe_read_req => zeropad_input_pipe_pipe_read_req(0 downto 0),
      zeropad_input_pipe_pipe_read_ack => zeropad_input_pipe_pipe_read_ack(0 downto 0),
      zeropad_input_pipe_pipe_read_data => zeropad_input_pipe_pipe_read_data(7 downto 0),
      zeropad_output_pipe_pipe_write_req => zeropad_output_pipe_pipe_write_req(0 downto 0),
      zeropad_output_pipe_pipe_write_ack => zeropad_output_pipe_pipe_write_ack(0 downto 0),
      zeropad_output_pipe_pipe_write_data => zeropad_output_pipe_pipe_write_data(7 downto 0),
      sendOutput_call_reqs => sendOutput_call_reqs(0 downto 0),
      sendOutput_call_acks => sendOutput_call_acks(0 downto 0),
      sendOutput_call_data => sendOutput_call_data(31 downto 0),
      sendOutput_call_tag => sendOutput_call_tag(0 downto 0),
      sendOutput_return_reqs => sendOutput_return_reqs(0 downto 0),
      sendOutput_return_acks => sendOutput_return_acks(0 downto 0),
      sendOutput_return_tag => sendOutput_return_tag(0 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      tag_in => zeropad3D_tag_in,
      tag_out => zeropad3D_tag_out-- 
    ); -- 
  -- module will be run forever 
  zeropad3D_tag_in <= (others => '0');
  zeropad3D_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => zeropad3D_start_req, start_ack => zeropad3D_start_ack,  fin_req => zeropad3D_fin_req,  fin_ack => zeropad3D_fin_ack);
  zeropad_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe zeropad_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => zeropad_input_pipe_pipe_read_req,
      read_ack => zeropad_input_pipe_pipe_read_ack,
      read_data => zeropad_input_pipe_pipe_read_data,
      write_req => zeropad_input_pipe_pipe_write_req,
      write_ack => zeropad_input_pipe_pipe_write_ack,
      write_data => zeropad_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  zeropad_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe zeropad_output_pipe",
      num_reads => 1,
      num_writes => 2,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => zeropad_output_pipe_pipe_read_req,
      read_ack => zeropad_output_pipe_pipe_read_ack,
      read_data => zeropad_output_pipe_pipe_read_data,
      write_req => zeropad_output_pipe_pipe_write_req,
      write_ack => zeropad_output_pipe_pipe_write_ack,
      write_data => zeropad_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
