-- VHDL global package produced by vc2vhdl from virtual circuit (vc) description 
library ieee;
use ieee.std_logic_1164.all;
package ahir_system_global_package is -- 
  constant global_time_val_base_address : std_logic_vector(4 downto 0) := "00000";
  -- 
end package ahir_system_global_package;
