-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTranspose is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(10 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTranspose;
architecture convTranspose_arch of convTranspose is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTranspose_CP_39_start: Boolean;
  signal convTranspose_CP_39_symbol: Boolean;
  -- volatile/operator module components. 
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal WPIPE_Block1_start_1018_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1039_inst_req_1 : boolean;
  signal type_cast_728_inst_req_0 : boolean;
  signal type_cast_728_inst_req_1 : boolean;
  signal type_cast_728_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_742_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1095_inst_ack_1 : boolean;
  signal type_cast_575_inst_ack_1 : boolean;
  signal type_cast_728_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1059_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1009_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1039_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_589_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_589_inst_req_1 : boolean;
  signal type_cast_521_inst_ack_1 : boolean;
  signal type_cast_575_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_724_inst_req_0 : boolean;
  signal array_obj_ref_689_index_offset_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_742_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_589_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_589_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_535_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_535_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_535_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_535_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_35_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1006_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_35_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_35_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_35_inst_ack_1 : boolean;
  signal array_obj_ref_689_index_offset_req_1 : boolean;
  signal type_cast_39_inst_req_0 : boolean;
  signal type_cast_39_inst_ack_0 : boolean;
  signal type_cast_39_inst_req_1 : boolean;
  signal type_cast_39_inst_ack_1 : boolean;
  signal addr_of_690_final_reg_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_135_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_135_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_571_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_135_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_135_inst_ack_1 : boolean;
  signal type_cast_710_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_48_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_48_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_48_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_48_inst_ack_1 : boolean;
  signal type_cast_710_inst_ack_1 : boolean;
  signal type_cast_660_inst_ack_0 : boolean;
  signal type_cast_52_inst_req_0 : boolean;
  signal type_cast_52_inst_ack_0 : boolean;
  signal type_cast_52_inst_req_1 : boolean;
  signal type_cast_52_inst_ack_1 : boolean;
  signal type_cast_575_inst_ack_0 : boolean;
  signal type_cast_1283_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1018_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_60_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1071_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_60_inst_ack_0 : boolean;
  signal type_cast_575_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_60_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_60_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_706_inst_ack_0 : boolean;
  signal type_cast_1050_inst_ack_0 : boolean;
  signal type_cast_64_inst_req_0 : boolean;
  signal type_cast_64_inst_ack_0 : boolean;
  signal type_cast_64_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1071_inst_ack_0 : boolean;
  signal type_cast_64_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_73_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_73_inst_ack_0 : boolean;
  signal addr_of_690_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_73_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_73_inst_ack_1 : boolean;
  signal type_cast_710_inst_req_1 : boolean;
  signal type_cast_697_inst_ack_1 : boolean;
  signal type_cast_697_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_706_inst_req_0 : boolean;
  signal type_cast_660_inst_req_0 : boolean;
  signal type_cast_77_inst_req_0 : boolean;
  signal type_cast_77_inst_ack_0 : boolean;
  signal type_cast_77_inst_req_1 : boolean;
  signal type_cast_77_inst_ack_1 : boolean;
  signal addr_of_690_final_reg_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_85_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_85_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_85_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_85_inst_ack_1 : boolean;
  signal type_cast_697_inst_ack_0 : boolean;
  signal array_obj_ref_689_index_offset_ack_0 : boolean;
  signal WPIPE_Block0_start_1006_inst_req_0 : boolean;
  signal type_cast_89_inst_req_0 : boolean;
  signal type_cast_89_inst_ack_0 : boolean;
  signal type_cast_89_inst_req_1 : boolean;
  signal type_cast_89_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1303_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_98_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_98_inst_ack_0 : boolean;
  signal if_stmt_633_branch_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_98_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_98_inst_ack_1 : boolean;
  signal type_cast_697_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1006_inst_ack_0 : boolean;
  signal type_cast_1050_inst_req_1 : boolean;
  signal type_cast_102_inst_req_0 : boolean;
  signal type_cast_102_inst_ack_0 : boolean;
  signal type_cast_102_inst_req_1 : boolean;
  signal type_cast_102_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_724_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_110_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_110_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_571_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_110_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_110_inst_ack_1 : boolean;
  signal array_obj_ref_689_index_offset_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_607_inst_ack_1 : boolean;
  signal type_cast_114_inst_req_0 : boolean;
  signal type_cast_114_inst_ack_0 : boolean;
  signal type_cast_114_inst_req_1 : boolean;
  signal type_cast_114_inst_ack_1 : boolean;
  signal type_cast_1425_inst_ack_1 : boolean;
  signal type_cast_1425_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_724_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_571_inst_req_1 : boolean;
  signal if_stmt_633_branch_ack_1 : boolean;
  signal addr_of_690_final_reg_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_123_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_123_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_123_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_123_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1059_inst_ack_0 : boolean;
  signal type_cast_1050_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_607_inst_req_1 : boolean;
  signal type_cast_127_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1071_inst_req_1 : boolean;
  signal type_cast_127_inst_ack_0 : boolean;
  signal type_cast_127_inst_req_1 : boolean;
  signal type_cast_127_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_706_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1052_inst_req_0 : boolean;
  signal type_cast_340_inst_req_0 : boolean;
  signal type_cast_340_inst_ack_0 : boolean;
  signal type_cast_340_inst_req_1 : boolean;
  signal type_cast_340_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1009_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1021_inst_ack_1 : boolean;
  signal type_cast_1395_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_349_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_349_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1052_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_349_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_349_inst_ack_1 : boolean;
  signal type_cast_139_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1071_inst_ack_1 : boolean;
  signal type_cast_139_inst_ack_0 : boolean;
  signal type_cast_139_inst_req_1 : boolean;
  signal type_cast_139_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_706_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_571_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1027_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_148_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_148_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_148_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_148_inst_ack_1 : boolean;
  signal type_cast_710_inst_req_0 : boolean;
  signal type_cast_660_inst_ack_1 : boolean;
  signal type_cast_152_inst_req_0 : boolean;
  signal type_cast_152_inst_ack_0 : boolean;
  signal type_cast_152_inst_req_1 : boolean;
  signal type_cast_152_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_724_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_160_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_160_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_160_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_160_inst_ack_1 : boolean;
  signal type_cast_1050_inst_req_0 : boolean;
  signal type_cast_164_inst_req_0 : boolean;
  signal type_cast_164_inst_ack_0 : boolean;
  signal type_cast_164_inst_req_1 : boolean;
  signal type_cast_164_inst_ack_1 : boolean;
  signal if_stmt_633_branch_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_173_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_173_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_173_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_173_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_693_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1303_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_607_inst_ack_0 : boolean;
  signal type_cast_660_inst_req_1 : boolean;
  signal type_cast_177_inst_req_0 : boolean;
  signal type_cast_177_inst_ack_0 : boolean;
  signal type_cast_177_inst_req_1 : boolean;
  signal type_cast_177_inst_ack_1 : boolean;
  signal type_cast_557_inst_ack_1 : boolean;
  signal type_cast_557_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_185_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_185_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_185_inst_req_1 : boolean;
  signal WPIPE_Block0_start_1006_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_185_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_693_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_607_inst_req_0 : boolean;
  signal type_cast_189_inst_req_0 : boolean;
  signal type_cast_189_inst_ack_0 : boolean;
  signal type_cast_189_inst_req_1 : boolean;
  signal type_cast_189_inst_ack_1 : boolean;
  signal type_cast_557_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1027_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_198_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_198_inst_ack_0 : boolean;
  signal type_cast_557_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_198_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_198_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1059_inst_req_1 : boolean;
  signal type_cast_202_inst_req_0 : boolean;
  signal type_cast_202_inst_ack_0 : boolean;
  signal type_cast_202_inst_req_1 : boolean;
  signal type_cast_202_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1021_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1027_inst_ack_0 : boolean;
  signal type_cast_211_inst_req_0 : boolean;
  signal type_cast_211_inst_ack_0 : boolean;
  signal type_cast_521_inst_req_1 : boolean;
  signal type_cast_211_inst_req_1 : boolean;
  signal type_cast_211_inst_ack_1 : boolean;
  signal ptr_deref_619_store_0_ack_1 : boolean;
  signal type_cast_215_inst_req_0 : boolean;
  signal type_cast_215_inst_ack_0 : boolean;
  signal type_cast_215_inst_req_1 : boolean;
  signal type_cast_215_inst_ack_1 : boolean;
  signal ptr_deref_619_store_0_req_1 : boolean;
  signal WPIPE_Block1_start_1059_inst_ack_1 : boolean;
  signal type_cast_219_inst_req_0 : boolean;
  signal type_cast_219_inst_ack_0 : boolean;
  signal type_cast_219_inst_req_1 : boolean;
  signal type_cast_219_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_553_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_553_inst_req_1 : boolean;
  signal type_cast_256_inst_req_0 : boolean;
  signal type_cast_256_inst_ack_0 : boolean;
  signal type_cast_256_inst_req_1 : boolean;
  signal type_cast_256_inst_ack_1 : boolean;
  signal type_cast_593_inst_ack_1 : boolean;
  signal type_cast_593_inst_req_1 : boolean;
  signal type_cast_260_inst_req_0 : boolean;
  signal type_cast_260_inst_ack_0 : boolean;
  signal type_cast_521_inst_ack_0 : boolean;
  signal type_cast_260_inst_req_1 : boolean;
  signal type_cast_260_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_553_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_553_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1080_inst_req_0 : boolean;
  signal type_cast_264_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1074_inst_req_0 : boolean;
  signal type_cast_264_inst_ack_0 : boolean;
  signal type_cast_521_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1009_inst_ack_1 : boolean;
  signal type_cast_264_inst_req_1 : boolean;
  signal type_cast_264_inst_ack_1 : boolean;
  signal type_cast_593_inst_ack_0 : boolean;
  signal type_cast_593_inst_req_0 : boolean;
  signal type_cast_268_inst_req_0 : boolean;
  signal type_cast_268_inst_ack_0 : boolean;
  signal type_cast_268_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1074_inst_ack_0 : boolean;
  signal type_cast_268_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1062_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_693_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_286_inst_req_0 : boolean;
  signal type_cast_611_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_286_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_286_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_286_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_693_inst_req_0 : boolean;
  signal type_cast_290_inst_req_0 : boolean;
  signal type_cast_611_inst_req_1 : boolean;
  signal type_cast_290_inst_ack_0 : boolean;
  signal type_cast_290_inst_req_1 : boolean;
  signal type_cast_290_inst_ack_1 : boolean;
  signal type_cast_539_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_299_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_299_inst_ack_0 : boolean;
  signal type_cast_539_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_299_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_299_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1080_inst_ack_0 : boolean;
  signal type_cast_303_inst_req_0 : boolean;
  signal type_cast_303_inst_ack_0 : boolean;
  signal type_cast_303_inst_req_1 : boolean;
  signal type_cast_611_inst_ack_0 : boolean;
  signal type_cast_303_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_311_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_311_inst_ack_0 : boolean;
  signal type_cast_539_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_311_inst_req_1 : boolean;
  signal type_cast_611_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_311_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1021_inst_ack_0 : boolean;
  signal type_cast_315_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1074_inst_req_1 : boolean;
  signal type_cast_315_inst_ack_0 : boolean;
  signal type_cast_315_inst_req_1 : boolean;
  signal type_cast_315_inst_ack_1 : boolean;
  signal type_cast_539_inst_req_0 : boolean;
  signal ptr_deref_619_store_0_ack_0 : boolean;
  signal ptr_deref_619_store_0_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_324_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_324_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_324_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1074_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_324_inst_ack_1 : boolean;
  signal type_cast_328_inst_req_0 : boolean;
  signal type_cast_328_inst_ack_0 : boolean;
  signal type_cast_328_inst_req_1 : boolean;
  signal type_cast_328_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1083_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_336_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_336_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_336_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_336_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1009_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1021_inst_req_1 : boolean;
  signal WPIPE_Block0_start_1012_inst_req_0 : boolean;
  signal type_cast_353_inst_req_0 : boolean;
  signal type_cast_353_inst_ack_0 : boolean;
  signal type_cast_353_inst_req_1 : boolean;
  signal type_cast_353_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1083_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_361_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_361_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_361_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_361_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1052_inst_req_1 : boolean;
  signal type_cast_365_inst_req_0 : boolean;
  signal type_cast_365_inst_ack_0 : boolean;
  signal addr_of_1367_final_reg_req_0 : boolean;
  signal type_cast_365_inst_req_1 : boolean;
  signal type_cast_365_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1024_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1052_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_374_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_374_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1024_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_374_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_374_inst_ack_1 : boolean;
  signal type_cast_378_inst_req_0 : boolean;
  signal type_cast_378_inst_ack_0 : boolean;
  signal type_cast_378_inst_req_1 : boolean;
  signal type_cast_378_inst_ack_1 : boolean;
  signal type_cast_1425_inst_req_0 : boolean;
  signal type_cast_1395_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_386_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_386_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_386_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_386_inst_ack_1 : boolean;
  signal type_cast_390_inst_req_0 : boolean;
  signal type_cast_390_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1012_inst_ack_0 : boolean;
  signal type_cast_390_inst_req_1 : boolean;
  signal type_cast_390_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1083_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_399_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_399_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_399_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_399_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1024_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1024_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1080_inst_req_1 : boolean;
  signal type_cast_1057_inst_req_0 : boolean;
  signal type_cast_403_inst_req_0 : boolean;
  signal type_cast_403_inst_ack_0 : boolean;
  signal type_cast_403_inst_req_1 : boolean;
  signal type_cast_1375_inst_ack_0 : boolean;
  signal type_cast_403_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1092_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1080_inst_ack_1 : boolean;
  signal type_cast_1425_inst_req_1 : boolean;
  signal type_cast_1057_inst_ack_0 : boolean;
  signal if_stmt_417_branch_req_0 : boolean;
  signal if_stmt_417_branch_ack_1 : boolean;
  signal if_stmt_417_branch_ack_0 : boolean;
  signal if_stmt_432_branch_req_0 : boolean;
  signal if_stmt_432_branch_ack_1 : boolean;
  signal if_stmt_432_branch_ack_0 : boolean;
  signal type_cast_453_inst_req_0 : boolean;
  signal type_cast_453_inst_ack_0 : boolean;
  signal type_cast_453_inst_req_1 : boolean;
  signal type_cast_453_inst_ack_1 : boolean;
  signal array_obj_ref_482_index_offset_req_0 : boolean;
  signal array_obj_ref_482_index_offset_ack_0 : boolean;
  signal array_obj_ref_482_index_offset_req_1 : boolean;
  signal array_obj_ref_482_index_offset_ack_1 : boolean;
  signal addr_of_483_final_reg_req_0 : boolean;
  signal addr_of_483_final_reg_ack_0 : boolean;
  signal addr_of_483_final_reg_req_1 : boolean;
  signal addr_of_483_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_486_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_486_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_486_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_486_inst_ack_1 : boolean;
  signal type_cast_490_inst_req_0 : boolean;
  signal type_cast_490_inst_ack_0 : boolean;
  signal type_cast_490_inst_req_1 : boolean;
  signal type_cast_490_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_499_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_499_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_499_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_499_inst_ack_1 : boolean;
  signal type_cast_503_inst_req_0 : boolean;
  signal type_cast_503_inst_ack_0 : boolean;
  signal type_cast_503_inst_req_1 : boolean;
  signal type_cast_503_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_517_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_517_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_517_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_517_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_742_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_742_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1039_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1039_inst_req_0 : boolean;
  signal type_cast_746_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1068_inst_ack_1 : boolean;
  signal type_cast_746_inst_ack_0 : boolean;
  signal type_cast_746_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1068_inst_req_1 : boolean;
  signal type_cast_746_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1095_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1092_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1018_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1095_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_760_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_760_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1018_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_760_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_760_inst_ack_1 : boolean;
  signal type_cast_1375_inst_req_0 : boolean;
  signal type_cast_764_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1068_inst_ack_0 : boolean;
  signal type_cast_764_inst_ack_0 : boolean;
  signal type_cast_764_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1068_inst_req_0 : boolean;
  signal type_cast_764_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1095_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1092_inst_req_1 : boolean;
  signal type_cast_1395_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_778_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_778_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_778_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_778_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1089_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1089_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1036_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1086_inst_ack_1 : boolean;
  signal type_cast_782_inst_req_0 : boolean;
  signal type_cast_782_inst_ack_0 : boolean;
  signal type_cast_782_inst_req_1 : boolean;
  signal type_cast_782_inst_ack_1 : boolean;
  signal addr_of_1367_final_reg_ack_0 : boolean;
  signal WPIPE_Block1_start_1036_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_796_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_796_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_796_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_796_inst_ack_1 : boolean;
  signal type_cast_1283_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1089_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1036_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1036_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1089_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1086_inst_req_1 : boolean;
  signal type_cast_800_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1065_inst_ack_1 : boolean;
  signal type_cast_800_inst_ack_0 : boolean;
  signal type_cast_800_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1065_inst_req_1 : boolean;
  signal type_cast_800_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1077_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_814_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_814_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1015_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_814_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_814_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1015_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1077_inst_req_1 : boolean;
  signal type_cast_818_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1065_inst_ack_0 : boolean;
  signal type_cast_818_inst_ack_0 : boolean;
  signal type_cast_818_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1065_inst_req_0 : boolean;
  signal type_cast_818_inst_ack_1 : boolean;
  signal type_cast_1395_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1092_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1300_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1077_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1077_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1033_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1033_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1027_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1086_inst_ack_0 : boolean;
  signal ptr_deref_826_store_0_req_0 : boolean;
  signal ptr_deref_826_store_0_ack_0 : boolean;
  signal WPIPE_Block0_start_1002_inst_ack_1 : boolean;
  signal ptr_deref_826_store_0_req_1 : boolean;
  signal WPIPE_Block1_start_1033_inst_ack_0 : boolean;
  signal ptr_deref_826_store_0_ack_1 : boolean;
  signal WPIPE_Block0_start_1002_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1033_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1015_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1083_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1030_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1015_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1086_inst_req_0 : boolean;
  signal if_stmt_840_branch_req_0 : boolean;
  signal WPIPE_Block1_start_1030_inst_req_1 : boolean;
  signal if_stmt_840_branch_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1288_inst_ack_0 : boolean;
  signal if_stmt_840_branch_ack_0 : boolean;
  signal type_cast_851_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1062_inst_ack_1 : boolean;
  signal type_cast_851_inst_ack_0 : boolean;
  signal type_cast_851_inst_req_1 : boolean;
  signal type_cast_851_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1300_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1030_inst_ack_0 : boolean;
  signal type_cast_855_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1062_inst_req_1 : boolean;
  signal type_cast_855_inst_ack_0 : boolean;
  signal type_cast_855_inst_req_1 : boolean;
  signal type_cast_855_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1030_inst_req_0 : boolean;
  signal type_cast_859_inst_req_0 : boolean;
  signal type_cast_859_inst_ack_0 : boolean;
  signal type_cast_859_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1062_inst_ack_0 : boolean;
  signal type_cast_859_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1012_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1012_inst_req_1 : boolean;
  signal type_cast_1057_inst_ack_1 : boolean;
  signal if_stmt_877_branch_req_0 : boolean;
  signal type_cast_1057_inst_req_1 : boolean;
  signal if_stmt_877_branch_ack_1 : boolean;
  signal if_stmt_877_branch_ack_0 : boolean;
  signal type_cast_1283_inst_ack_1 : boolean;
  signal type_cast_904_inst_req_0 : boolean;
  signal type_cast_904_inst_ack_0 : boolean;
  signal type_cast_904_inst_req_1 : boolean;
  signal type_cast_904_inst_ack_1 : boolean;
  signal type_cast_1375_inst_req_1 : boolean;
  signal type_cast_1405_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1300_inst_req_1 : boolean;
  signal array_obj_ref_933_index_offset_req_0 : boolean;
  signal array_obj_ref_933_index_offset_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1300_inst_ack_1 : boolean;
  signal array_obj_ref_933_index_offset_req_1 : boolean;
  signal array_obj_ref_933_index_offset_ack_1 : boolean;
  signal array_obj_ref_1366_index_offset_req_0 : boolean;
  signal type_cast_1375_inst_ack_1 : boolean;
  signal addr_of_934_final_reg_req_0 : boolean;
  signal addr_of_934_final_reg_ack_0 : boolean;
  signal addr_of_934_final_reg_req_1 : boolean;
  signal addr_of_934_final_reg_ack_1 : boolean;
  signal type_cast_1405_inst_ack_0 : boolean;
  signal array_obj_ref_1366_index_offset_ack_0 : boolean;
  signal array_obj_ref_1366_index_offset_req_1 : boolean;
  signal addr_of_1367_final_reg_req_1 : boolean;
  signal array_obj_ref_1366_index_offset_ack_1 : boolean;
  signal ptr_deref_937_store_0_req_0 : boolean;
  signal ptr_deref_937_store_0_ack_0 : boolean;
  signal ptr_deref_937_store_0_req_1 : boolean;
  signal ptr_deref_937_store_0_ack_1 : boolean;
  signal addr_of_1367_final_reg_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1288_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1288_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1285_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1285_inst_ack_0 : boolean;
  signal if_stmt_952_branch_req_0 : boolean;
  signal if_stmt_952_branch_ack_1 : boolean;
  signal if_stmt_952_branch_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1303_inst_req_0 : boolean;
  signal call_stmt_963_call_req_0 : boolean;
  signal call_stmt_963_call_ack_0 : boolean;
  signal type_cast_1445_inst_req_0 : boolean;
  signal call_stmt_963_call_req_1 : boolean;
  signal call_stmt_963_call_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1303_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1285_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1285_inst_ack_1 : boolean;
  signal type_cast_968_inst_req_0 : boolean;
  signal type_cast_968_inst_ack_0 : boolean;
  signal type_cast_968_inst_req_1 : boolean;
  signal type_cast_968_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_971_inst_req_0 : boolean;
  signal WPIPE_Block0_start_971_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_971_inst_req_1 : boolean;
  signal WPIPE_Block0_start_971_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_974_inst_req_0 : boolean;
  signal WPIPE_Block0_start_974_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_974_inst_req_1 : boolean;
  signal WPIPE_Block0_start_974_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_977_inst_req_0 : boolean;
  signal WPIPE_Block0_start_977_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_977_inst_req_1 : boolean;
  signal WPIPE_Block0_start_977_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_980_inst_req_0 : boolean;
  signal WPIPE_Block0_start_980_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_980_inst_req_1 : boolean;
  signal WPIPE_Block0_start_980_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_983_inst_req_0 : boolean;
  signal WPIPE_Block0_start_983_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_983_inst_req_1 : boolean;
  signal WPIPE_Block0_start_983_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_986_inst_req_0 : boolean;
  signal WPIPE_Block0_start_986_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_986_inst_req_1 : boolean;
  signal WPIPE_Block0_start_986_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_989_inst_req_0 : boolean;
  signal WPIPE_Block0_start_989_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_989_inst_req_1 : boolean;
  signal WPIPE_Block0_start_989_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_992_inst_req_0 : boolean;
  signal WPIPE_Block0_start_992_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_992_inst_req_1 : boolean;
  signal WPIPE_Block0_start_992_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_995_inst_req_0 : boolean;
  signal WPIPE_Block0_start_995_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_995_inst_req_1 : boolean;
  signal WPIPE_Block0_start_995_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_998_inst_req_0 : boolean;
  signal WPIPE_Block0_start_998_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_998_inst_req_1 : boolean;
  signal WPIPE_Block0_start_998_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1002_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1002_inst_ack_0 : boolean;
  signal type_cast_1106_inst_req_0 : boolean;
  signal type_cast_1106_inst_ack_0 : boolean;
  signal type_cast_1106_inst_req_1 : boolean;
  signal type_cast_1106_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1108_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1108_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1108_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1108_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1450_inst_ack_1 : boolean;
  signal type_cast_1435_inst_ack_1 : boolean;
  signal type_cast_1113_inst_req_0 : boolean;
  signal type_cast_1113_inst_ack_0 : boolean;
  signal type_cast_1435_inst_req_1 : boolean;
  signal type_cast_1113_inst_req_1 : boolean;
  signal type_cast_1113_inst_ack_1 : boolean;
  signal type_cast_1385_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1115_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1115_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1288_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1115_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1115_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1450_inst_req_1 : boolean;
  signal type_cast_1385_inst_req_1 : boolean;
  signal type_cast_1337_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1118_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1118_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1297_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1118_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1118_inst_ack_1 : boolean;
  signal type_cast_1337_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1121_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1121_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1297_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1121_inst_req_1 : boolean;
  signal ptr_deref_1371_load_0_ack_1 : boolean;
  signal WPIPE_Block2_start_1121_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1450_inst_ack_0 : boolean;
  signal type_cast_1385_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1124_inst_req_0 : boolean;
  signal ptr_deref_1371_load_0_req_1 : boolean;
  signal WPIPE_Block2_start_1124_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1124_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1124_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1450_inst_req_0 : boolean;
  signal type_cast_1385_inst_req_0 : boolean;
  signal type_cast_1415_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1127_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1127_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1127_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1127_inst_ack_1 : boolean;
  signal type_cast_1337_inst_ack_0 : boolean;
  signal type_cast_1415_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1130_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1130_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1297_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1130_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1130_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1297_inst_req_0 : boolean;
  signal type_cast_1337_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1133_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1133_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1133_inst_req_1 : boolean;
  signal ptr_deref_1371_load_0_ack_0 : boolean;
  signal WPIPE_Block3_start_1133_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1453_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1136_inst_req_0 : boolean;
  signal ptr_deref_1371_load_0_req_0 : boolean;
  signal WPIPE_Block3_start_1136_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1136_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1136_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1453_inst_req_1 : boolean;
  signal type_cast_1415_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1139_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1139_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1139_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1139_inst_ack_1 : boolean;
  signal type_cast_1415_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1142_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1142_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1294_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1142_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1142_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1294_inst_req_1 : boolean;
  signal if_stmt_1310_branch_ack_0 : boolean;
  signal WPIPE_Block3_start_1145_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1145_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1145_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1145_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1447_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1447_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1148_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1148_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1294_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1148_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1148_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1294_inst_req_0 : boolean;
  signal if_stmt_1310_branch_ack_1 : boolean;
  signal WPIPE_Block3_start_1151_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1151_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1151_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1151_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1447_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1447_inst_req_0 : boolean;
  signal if_stmt_1310_branch_req_0 : boolean;
  signal type_cast_1162_inst_req_0 : boolean;
  signal type_cast_1162_inst_ack_0 : boolean;
  signal type_cast_1435_inst_ack_0 : boolean;
  signal type_cast_1162_inst_req_1 : boolean;
  signal type_cast_1162_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1164_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1164_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1164_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1164_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1453_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1306_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1306_inst_req_1 : boolean;
  signal type_cast_1435_inst_req_0 : boolean;
  signal type_cast_1169_inst_req_0 : boolean;
  signal type_cast_1169_inst_ack_0 : boolean;
  signal type_cast_1169_inst_req_1 : boolean;
  signal type_cast_1169_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1291_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1291_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1171_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1171_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1171_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1171_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1453_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1306_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1174_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1174_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1291_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1174_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1174_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1291_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1306_inst_req_0 : boolean;
  signal type_cast_1405_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1177_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1177_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1177_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1177_inst_ack_1 : boolean;
  signal type_cast_1445_inst_ack_1 : boolean;
  signal type_cast_1445_inst_req_1 : boolean;
  signal type_cast_1405_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1180_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1180_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1180_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1180_inst_ack_1 : boolean;
  signal type_cast_1445_inst_ack_0 : boolean;
  signal RPIPE_Block0_done_1184_inst_req_0 : boolean;
  signal RPIPE_Block0_done_1184_inst_ack_0 : boolean;
  signal RPIPE_Block0_done_1184_inst_req_1 : boolean;
  signal RPIPE_Block0_done_1184_inst_ack_1 : boolean;
  signal RPIPE_Block1_done_1187_inst_req_0 : boolean;
  signal RPIPE_Block1_done_1187_inst_ack_0 : boolean;
  signal RPIPE_Block1_done_1187_inst_req_1 : boolean;
  signal RPIPE_Block1_done_1187_inst_ack_1 : boolean;
  signal RPIPE_Block2_done_1190_inst_req_0 : boolean;
  signal RPIPE_Block2_done_1190_inst_ack_0 : boolean;
  signal RPIPE_Block2_done_1190_inst_req_1 : boolean;
  signal RPIPE_Block2_done_1190_inst_ack_1 : boolean;
  signal RPIPE_Block3_done_1193_inst_req_0 : boolean;
  signal RPIPE_Block3_done_1193_inst_ack_0 : boolean;
  signal RPIPE_Block3_done_1193_inst_req_1 : boolean;
  signal RPIPE_Block3_done_1193_inst_ack_1 : boolean;
  signal call_stmt_1197_call_req_0 : boolean;
  signal call_stmt_1197_call_ack_0 : boolean;
  signal call_stmt_1197_call_req_1 : boolean;
  signal call_stmt_1197_call_ack_1 : boolean;
  signal type_cast_1201_inst_req_0 : boolean;
  signal type_cast_1201_inst_ack_0 : boolean;
  signal type_cast_1201_inst_req_1 : boolean;
  signal type_cast_1201_inst_ack_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1208_inst_req_0 : boolean;
  signal WPIPE_elapsed_time_pipe_1208_inst_ack_0 : boolean;
  signal WPIPE_elapsed_time_pipe_1208_inst_req_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1208_inst_ack_1 : boolean;
  signal type_cast_1213_inst_req_0 : boolean;
  signal type_cast_1213_inst_ack_0 : boolean;
  signal type_cast_1213_inst_req_1 : boolean;
  signal type_cast_1213_inst_ack_1 : boolean;
  signal type_cast_1223_inst_req_0 : boolean;
  signal type_cast_1223_inst_ack_0 : boolean;
  signal type_cast_1223_inst_req_1 : boolean;
  signal type_cast_1223_inst_ack_1 : boolean;
  signal type_cast_1233_inst_req_0 : boolean;
  signal type_cast_1233_inst_ack_0 : boolean;
  signal type_cast_1233_inst_req_1 : boolean;
  signal type_cast_1233_inst_ack_1 : boolean;
  signal type_cast_1243_inst_req_0 : boolean;
  signal type_cast_1243_inst_ack_0 : boolean;
  signal type_cast_1243_inst_req_1 : boolean;
  signal type_cast_1243_inst_ack_1 : boolean;
  signal type_cast_1253_inst_req_0 : boolean;
  signal type_cast_1253_inst_ack_0 : boolean;
  signal type_cast_1253_inst_req_1 : boolean;
  signal type_cast_1253_inst_ack_1 : boolean;
  signal type_cast_1263_inst_req_0 : boolean;
  signal type_cast_1263_inst_ack_0 : boolean;
  signal type_cast_1263_inst_req_1 : boolean;
  signal type_cast_1263_inst_ack_1 : boolean;
  signal type_cast_1273_inst_req_0 : boolean;
  signal type_cast_1273_inst_ack_0 : boolean;
  signal type_cast_1273_inst_req_1 : boolean;
  signal type_cast_1273_inst_ack_1 : boolean;
  signal type_cast_1283_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1456_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1456_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1456_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1456_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1459_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1459_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1459_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1459_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1462_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1462_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1462_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1462_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1465_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1465_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1465_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1465_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1468_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1468_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1468_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1468_inst_ack_1 : boolean;
  signal if_stmt_1482_branch_req_0 : boolean;
  signal if_stmt_1482_branch_ack_1 : boolean;
  signal if_stmt_1482_branch_ack_0 : boolean;
  signal phi_stmt_470_req_0 : boolean;
  signal type_cast_476_inst_req_0 : boolean;
  signal type_cast_476_inst_ack_0 : boolean;
  signal type_cast_476_inst_req_1 : boolean;
  signal type_cast_476_inst_ack_1 : boolean;
  signal phi_stmt_470_req_1 : boolean;
  signal phi_stmt_470_ack_0 : boolean;
  signal phi_stmt_677_req_0 : boolean;
  signal type_cast_683_inst_req_0 : boolean;
  signal type_cast_683_inst_ack_0 : boolean;
  signal type_cast_683_inst_req_1 : boolean;
  signal type_cast_683_inst_ack_1 : boolean;
  signal phi_stmt_677_req_1 : boolean;
  signal phi_stmt_677_ack_0 : boolean;
  signal phi_stmt_921_req_1 : boolean;
  signal type_cast_924_inst_req_0 : boolean;
  signal type_cast_924_inst_ack_0 : boolean;
  signal type_cast_924_inst_req_1 : boolean;
  signal type_cast_924_inst_ack_1 : boolean;
  signal phi_stmt_921_req_0 : boolean;
  signal phi_stmt_921_ack_0 : boolean;
  signal phi_stmt_1354_req_0 : boolean;
  signal type_cast_1360_inst_req_0 : boolean;
  signal type_cast_1360_inst_ack_0 : boolean;
  signal type_cast_1360_inst_req_1 : boolean;
  signal type_cast_1360_inst_ack_1 : boolean;
  signal phi_stmt_1354_req_1 : boolean;
  signal phi_stmt_1354_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTranspose_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTranspose_CP_39_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTranspose_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_39_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTranspose_CP_39_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_39_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTranspose_CP_39: Block -- control-path 
    signal convTranspose_CP_39_elements: BooleanArray(499 downto 0);
    -- 
  begin -- 
    convTranspose_CP_39_elements(0) <= convTranspose_CP_39_start;
    convTranspose_CP_39_symbol <= convTranspose_CP_39_elements(499);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	52 
    -- CP-element group 0: 	40 
    -- CP-element group 0: 	48 
    -- CP-element group 0: 	44 
    -- CP-element group 0: 	56 
    -- CP-element group 0: 	59 
    -- CP-element group 0: 	62 
    -- CP-element group 0: 	65 
    -- CP-element group 0: 	68 
    -- CP-element group 0: 	71 
    -- CP-element group 0: 	74 
    -- CP-element group 0: 	77 
    -- CP-element group 0: 	81 
    -- CP-element group 0: 	85 
    -- CP-element group 0: 	89 
    -- CP-element group 0: 	93 
    -- CP-element group 0: 	97 
    -- CP-element group 0: 	101 
    -- CP-element group 0: 	105 
    -- CP-element group 0: 	109 
    -- CP-element group 0: 	113 
    -- CP-element group 0: 	117 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	12 
    -- CP-element group 0: 	16 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	24 
    -- CP-element group 0: 	28 
    -- CP-element group 0: 	32 
    -- CP-element group 0: 	36 
    -- CP-element group 0:  members (101) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_33/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/branch_block_stmt_33__entry__
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416__entry__
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_35_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_35_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_35_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_39_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_39_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_39_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_52_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_52_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_52_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_64_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_64_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_64_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_77_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_77_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_77_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_89_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_89_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_89_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_102_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_102_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_102_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_114_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_114_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_114_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_127_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_127_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_127_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_340_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_340_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_340_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_139_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_139_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_139_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_152_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_152_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_152_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_164_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_328_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_164_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_164_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_177_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_177_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_177_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_189_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_189_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_189_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_202_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_202_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_202_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_211_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_211_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_211_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_215_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_215_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_215_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_219_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_219_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_219_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_256_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_256_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_256_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_260_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_260_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_260_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_264_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_264_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_264_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_268_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_268_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_268_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_290_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_290_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_290_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_303_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_303_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_303_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_315_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_315_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_315_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_328_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_328_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_353_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_353_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_353_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_365_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_365_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_365_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_378_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_378_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_378_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_390_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_390_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_390_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_403_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_403_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_403_Update/cr
      -- 
    rr_135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => RPIPE_ConvTranspose_input_pipe_35_inst_req_0); -- 
    cr_154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_39_inst_req_1); -- 
    cr_182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_52_inst_req_1); -- 
    cr_210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_64_inst_req_1); -- 
    cr_238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_77_inst_req_1); -- 
    cr_266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_89_inst_req_1); -- 
    cr_294_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_294_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_102_inst_req_1); -- 
    cr_322_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_322_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_114_inst_req_1); -- 
    cr_350_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_350_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_127_inst_req_1); -- 
    cr_756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_340_inst_req_1); -- 
    cr_378_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_378_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_139_inst_req_1); -- 
    cr_406_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_406_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_152_inst_req_1); -- 
    cr_434_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_434_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_164_inst_req_1); -- 
    cr_462_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_462_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_177_inst_req_1); -- 
    cr_490_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_490_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_189_inst_req_1); -- 
    cr_518_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_518_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_202_inst_req_1); -- 
    cr_532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_211_inst_req_1); -- 
    cr_546_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_546_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_215_inst_req_1); -- 
    cr_560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_219_inst_req_1); -- 
    cr_574_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_574_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_256_inst_req_1); -- 
    cr_588_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_588_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_260_inst_req_1); -- 
    cr_602_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_602_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_264_inst_req_1); -- 
    cr_616_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_616_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_268_inst_req_1); -- 
    cr_644_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_644_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_290_inst_req_1); -- 
    cr_672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_303_inst_req_1); -- 
    cr_700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_315_inst_req_1); -- 
    cr_728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_328_inst_req_1); -- 
    cr_784_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_784_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_353_inst_req_1); -- 
    cr_812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_365_inst_req_1); -- 
    cr_840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_378_inst_req_1); -- 
    cr_868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_390_inst_req_1); -- 
    cr_896_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_896_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_403_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_35_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_35_update_start_
      -- CP-element group 1: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_35_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_35_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_35_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_35_Update/cr
      -- 
    ra_136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_35_inst_ack_0, ack => convTranspose_CP_39_elements(1)); -- 
    cr_140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(1), ack => RPIPE_ConvTranspose_input_pipe_35_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_48_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_48_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_35_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_35_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_35_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_39_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_39_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_39_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_48_Sample/rr
      -- 
    ca_141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_35_inst_ack_1, ack => convTranspose_CP_39_elements(2)); -- 
    rr_149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(2), ack => type_cast_39_inst_req_0); -- 
    rr_163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(2), ack => RPIPE_ConvTranspose_input_pipe_48_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_39_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_39_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_39_Sample/ra
      -- 
    ra_150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_39_inst_ack_0, ack => convTranspose_CP_39_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	57 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_39_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_39_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_39_Update/ca
      -- 
    ca_155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_39_inst_ack_1, ack => convTranspose_CP_39_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_48_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_48_update_start_
      -- CP-element group 5: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_48_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_48_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_48_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_48_Update/cr
      -- 
    ra_164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_48_inst_ack_0, ack => convTranspose_CP_39_elements(5)); -- 
    cr_168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(5), ack => RPIPE_ConvTranspose_input_pipe_48_inst_req_1); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_48_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_48_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_48_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_52_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_52_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_52_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_60_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_60_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_60_Sample/rr
      -- 
    ca_169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_48_inst_ack_1, ack => convTranspose_CP_39_elements(6)); -- 
    rr_177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(6), ack => type_cast_52_inst_req_0); -- 
    rr_191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(6), ack => RPIPE_ConvTranspose_input_pipe_60_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_52_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_52_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_52_Sample/ra
      -- 
    ra_178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_52_inst_ack_0, ack => convTranspose_CP_39_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	57 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_52_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_52_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_52_Update/ca
      -- 
    ca_183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_52_inst_ack_1, ack => convTranspose_CP_39_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_60_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_60_update_start_
      -- CP-element group 9: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_60_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_60_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_60_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_60_Update/cr
      -- 
    ra_192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_60_inst_ack_0, ack => convTranspose_CP_39_elements(9)); -- 
    cr_196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(9), ack => RPIPE_ConvTranspose_input_pipe_60_inst_req_1); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	13 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_60_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_60_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_60_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_64_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_64_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_64_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_73_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_73_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_73_Sample/rr
      -- 
    ca_197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_60_inst_ack_1, ack => convTranspose_CP_39_elements(10)); -- 
    rr_205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(10), ack => type_cast_64_inst_req_0); -- 
    rr_219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(10), ack => RPIPE_ConvTranspose_input_pipe_73_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_64_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_64_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_64_Sample/ra
      -- 
    ra_206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_64_inst_ack_0, ack => convTranspose_CP_39_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	60 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_64_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_64_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_64_Update/ca
      -- 
    ca_211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_64_inst_ack_1, ack => convTranspose_CP_39_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_73_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_73_update_start_
      -- CP-element group 13: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_73_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_73_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_73_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_73_Update/cr
      -- 
    ra_220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_73_inst_ack_0, ack => convTranspose_CP_39_elements(13)); -- 
    cr_224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(13), ack => RPIPE_ConvTranspose_input_pipe_73_inst_req_1); -- 
    -- CP-element group 14:  fork  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_73_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_73_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_73_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_77_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_77_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_77_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_85_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_85_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_85_Sample/rr
      -- 
    ca_225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_73_inst_ack_1, ack => convTranspose_CP_39_elements(14)); -- 
    rr_233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(14), ack => type_cast_77_inst_req_0); -- 
    rr_247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(14), ack => RPIPE_ConvTranspose_input_pipe_85_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_77_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_77_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_77_Sample/ra
      -- 
    ra_234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_77_inst_ack_0, ack => convTranspose_CP_39_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	0 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	60 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_77_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_77_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_77_Update/ca
      -- 
    ca_239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_77_inst_ack_1, ack => convTranspose_CP_39_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_85_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_85_update_start_
      -- CP-element group 17: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_85_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_85_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_85_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_85_Update/cr
      -- 
    ra_248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_85_inst_ack_0, ack => convTranspose_CP_39_elements(17)); -- 
    cr_252_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_252_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(17), ack => RPIPE_ConvTranspose_input_pipe_85_inst_req_1); -- 
    -- CP-element group 18:  fork  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18: 	21 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_85_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_85_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_85_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_89_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_89_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_89_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_98_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_98_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_98_Sample/rr
      -- 
    ca_253_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_85_inst_ack_1, ack => convTranspose_CP_39_elements(18)); -- 
    rr_261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(18), ack => type_cast_89_inst_req_0); -- 
    rr_275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(18), ack => RPIPE_ConvTranspose_input_pipe_98_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_89_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_89_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_89_Sample/ra
      -- 
    ra_262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_89_inst_ack_0, ack => convTranspose_CP_39_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	63 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_89_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_89_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_89_Update/ca
      -- 
    ca_267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_89_inst_ack_1, ack => convTranspose_CP_39_elements(20)); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_98_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_98_update_start_
      -- CP-element group 21: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_98_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_98_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_98_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_98_Update/cr
      -- 
    ra_276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_98_inst_ack_0, ack => convTranspose_CP_39_elements(21)); -- 
    cr_280_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_280_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(21), ack => RPIPE_ConvTranspose_input_pipe_98_inst_req_1); -- 
    -- CP-element group 22:  fork  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22: 	25 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_98_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_98_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_98_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_102_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_102_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_102_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_110_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_110_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_110_Sample/rr
      -- 
    ca_281_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_98_inst_ack_1, ack => convTranspose_CP_39_elements(22)); -- 
    rr_289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(22), ack => type_cast_102_inst_req_0); -- 
    rr_303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(22), ack => RPIPE_ConvTranspose_input_pipe_110_inst_req_0); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_102_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_102_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_102_Sample/ra
      -- 
    ra_290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_102_inst_ack_0, ack => convTranspose_CP_39_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	0 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	63 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_102_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_102_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_102_Update/ca
      -- 
    ca_295_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_102_inst_ack_1, ack => convTranspose_CP_39_elements(24)); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	22 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_110_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_110_update_start_
      -- CP-element group 25: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_110_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_110_Sample/ra
      -- CP-element group 25: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_110_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_110_Update/cr
      -- 
    ra_304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_110_inst_ack_0, ack => convTranspose_CP_39_elements(25)); -- 
    cr_308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(25), ack => RPIPE_ConvTranspose_input_pipe_110_inst_req_1); -- 
    -- CP-element group 26:  fork  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: 	29 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_110_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_110_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_110_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_114_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_114_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_114_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_123_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_123_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_123_Sample/rr
      -- 
    ca_309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_110_inst_ack_1, ack => convTranspose_CP_39_elements(26)); -- 
    rr_317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(26), ack => type_cast_114_inst_req_0); -- 
    rr_331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(26), ack => RPIPE_ConvTranspose_input_pipe_123_inst_req_0); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_114_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_114_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_114_Sample/ra
      -- 
    ra_318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_114_inst_ack_0, ack => convTranspose_CP_39_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	0 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	66 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_114_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_114_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_114_Update/ca
      -- 
    ca_323_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_114_inst_ack_1, ack => convTranspose_CP_39_elements(28)); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	26 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_123_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_123_update_start_
      -- CP-element group 29: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_123_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_123_Sample/ra
      -- CP-element group 29: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_123_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_123_Update/cr
      -- 
    ra_332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_123_inst_ack_0, ack => convTranspose_CP_39_elements(29)); -- 
    cr_336_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_336_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(29), ack => RPIPE_ConvTranspose_input_pipe_123_inst_req_1); -- 
    -- CP-element group 30:  fork  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: 	33 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_135_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_135_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_123_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_123_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_123_Update/ca
      -- CP-element group 30: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_127_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_127_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_127_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_135_sample_start_
      -- 
    ca_337_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_123_inst_ack_1, ack => convTranspose_CP_39_elements(30)); -- 
    rr_345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(30), ack => type_cast_127_inst_req_0); -- 
    rr_359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(30), ack => RPIPE_ConvTranspose_input_pipe_135_inst_req_0); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_127_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_127_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_127_Sample/ra
      -- 
    ra_346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_127_inst_ack_0, ack => convTranspose_CP_39_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	0 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	66 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_127_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_127_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_127_Update/ca
      -- 
    ca_351_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_127_inst_ack_1, ack => convTranspose_CP_39_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	30 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_135_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_135_Sample/ra
      -- CP-element group 33: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_135_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_135_Update/cr
      -- CP-element group 33: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_135_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_135_update_start_
      -- 
    ra_360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_135_inst_ack_0, ack => convTranspose_CP_39_elements(33)); -- 
    cr_364_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_364_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(33), ack => RPIPE_ConvTranspose_input_pipe_135_inst_req_1); -- 
    -- CP-element group 34:  fork  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	37 
    -- CP-element group 34:  members (9) 
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_135_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_135_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_135_Update/ca
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_139_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_139_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_139_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_148_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_148_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_148_Sample/rr
      -- 
    ca_365_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_135_inst_ack_1, ack => convTranspose_CP_39_elements(34)); -- 
    rr_373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(34), ack => type_cast_139_inst_req_0); -- 
    rr_387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(34), ack => RPIPE_ConvTranspose_input_pipe_148_inst_req_0); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_139_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_139_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_139_Sample/ra
      -- 
    ra_374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_139_inst_ack_0, ack => convTranspose_CP_39_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	0 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	69 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_139_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_139_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_139_Update/ca
      -- 
    ca_379_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_139_inst_ack_1, ack => convTranspose_CP_39_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_148_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_148_update_start_
      -- CP-element group 37: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_148_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_148_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_148_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_148_Update/cr
      -- 
    ra_388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_148_inst_ack_0, ack => convTranspose_CP_39_elements(37)); -- 
    cr_392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(37), ack => RPIPE_ConvTranspose_input_pipe_148_inst_req_1); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	41 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_148_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_148_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_148_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_152_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_152_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_152_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_160_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_160_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_160_Sample/rr
      -- 
    ca_393_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_148_inst_ack_1, ack => convTranspose_CP_39_elements(38)); -- 
    rr_401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(38), ack => type_cast_152_inst_req_0); -- 
    rr_415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(38), ack => RPIPE_ConvTranspose_input_pipe_160_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_152_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_152_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_152_Sample/ra
      -- 
    ra_402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_152_inst_ack_0, ack => convTranspose_CP_39_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	0 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	69 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_152_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_152_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_152_Update/ca
      -- 
    ca_407_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_152_inst_ack_1, ack => convTranspose_CP_39_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	38 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_160_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_160_update_start_
      -- CP-element group 41: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_160_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_160_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_160_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_160_Update/cr
      -- 
    ra_416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_160_inst_ack_0, ack => convTranspose_CP_39_elements(41)); -- 
    cr_420_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_420_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(41), ack => RPIPE_ConvTranspose_input_pipe_160_inst_req_1); -- 
    -- CP-element group 42:  fork  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42: 	45 
    -- CP-element group 42:  members (9) 
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_160_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_160_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_160_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_164_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_164_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_164_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_173_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_173_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_173_Sample/rr
      -- 
    ca_421_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_160_inst_ack_1, ack => convTranspose_CP_39_elements(42)); -- 
    rr_429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(42), ack => type_cast_164_inst_req_0); -- 
    rr_443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(42), ack => RPIPE_ConvTranspose_input_pipe_173_inst_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_164_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_164_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_164_Sample/ra
      -- 
    ra_430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_164_inst_ack_0, ack => convTranspose_CP_39_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	0 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	72 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_164_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_164_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_164_Update/ca
      -- 
    ca_435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_164_inst_ack_1, ack => convTranspose_CP_39_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	42 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_173_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_173_update_start_
      -- CP-element group 45: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_173_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_173_Sample/ra
      -- CP-element group 45: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_173_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_173_Update/cr
      -- 
    ra_444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_173_inst_ack_0, ack => convTranspose_CP_39_elements(45)); -- 
    cr_448_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_448_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(45), ack => RPIPE_ConvTranspose_input_pipe_173_inst_req_1); -- 
    -- CP-element group 46:  fork  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46: 	49 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_173_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_173_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_173_Update/ca
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_177_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_177_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_177_Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_185_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_185_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_185_Sample/rr
      -- 
    ca_449_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_173_inst_ack_1, ack => convTranspose_CP_39_elements(46)); -- 
    rr_457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(46), ack => type_cast_177_inst_req_0); -- 
    rr_471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(46), ack => RPIPE_ConvTranspose_input_pipe_185_inst_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_177_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_177_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_177_Sample/ra
      -- 
    ra_458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_177_inst_ack_0, ack => convTranspose_CP_39_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	0 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	72 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_177_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_177_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_177_Update/ca
      -- 
    ca_463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_177_inst_ack_1, ack => convTranspose_CP_39_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	46 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_185_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_185_update_start_
      -- CP-element group 49: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_185_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_185_Sample/ra
      -- CP-element group 49: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_185_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_185_Update/cr
      -- 
    ra_472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_185_inst_ack_0, ack => convTranspose_CP_39_elements(49)); -- 
    cr_476_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_476_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(49), ack => RPIPE_ConvTranspose_input_pipe_185_inst_req_1); -- 
    -- CP-element group 50:  fork  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	53 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_185_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_185_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_185_Update/ca
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_189_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_189_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_189_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_198_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_198_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_198_Sample/rr
      -- 
    ca_477_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_185_inst_ack_1, ack => convTranspose_CP_39_elements(50)); -- 
    rr_485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(50), ack => type_cast_189_inst_req_0); -- 
    rr_499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(50), ack => RPIPE_ConvTranspose_input_pipe_198_inst_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_189_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_189_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_189_Sample/ra
      -- 
    ra_486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_189_inst_ack_0, ack => convTranspose_CP_39_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	0 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	75 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_189_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_189_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_189_Update/ca
      -- 
    ca_491_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_189_inst_ack_1, ack => convTranspose_CP_39_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	50 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (6) 
      -- CP-element group 53: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_198_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_198_update_start_
      -- CP-element group 53: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_198_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_198_Sample/ra
      -- CP-element group 53: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_198_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_198_Update/cr
      -- 
    ra_500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_198_inst_ack_0, ack => convTranspose_CP_39_elements(53)); -- 
    cr_504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(53), ack => RPIPE_ConvTranspose_input_pipe_198_inst_req_1); -- 
    -- CP-element group 54:  fork  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54: 	78 
    -- CP-element group 54:  members (9) 
      -- CP-element group 54: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_198_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_198_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_198_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_202_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_202_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_202_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_286_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_286_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_286_Sample/rr
      -- 
    ca_505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_198_inst_ack_1, ack => convTranspose_CP_39_elements(54)); -- 
    rr_513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(54), ack => type_cast_202_inst_req_0); -- 
    rr_625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(54), ack => RPIPE_ConvTranspose_input_pipe_286_inst_req_0); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_202_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_202_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_202_Sample/ra
      -- 
    ra_514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_202_inst_ack_0, ack => convTranspose_CP_39_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	0 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	75 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_202_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_202_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_202_Update/ca
      -- 
    ca_519_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_202_inst_ack_1, ack => convTranspose_CP_39_elements(56)); -- 
    -- CP-element group 57:  join  transition  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	4 
    -- CP-element group 57: 	8 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_211_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_211_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_211_Sample/rr
      -- 
    rr_527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(57), ack => type_cast_211_inst_req_0); -- 
    convTranspose_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(4) & convTranspose_CP_39_elements(8);
      gj_convTranspose_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_211_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_211_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_211_Sample/ra
      -- 
    ra_528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_211_inst_ack_0, ack => convTranspose_CP_39_elements(58)); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	0 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	118 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_211_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_211_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_211_Update/ca
      -- 
    ca_533_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_211_inst_ack_1, ack => convTranspose_CP_39_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	12 
    -- CP-element group 60: 	16 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_215_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_215_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_215_Sample/rr
      -- 
    rr_541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(60), ack => type_cast_215_inst_req_0); -- 
    convTranspose_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(12) & convTranspose_CP_39_elements(16);
      gj_convTranspose_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_215_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_215_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_215_Sample/ra
      -- 
    ra_542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_215_inst_ack_0, ack => convTranspose_CP_39_elements(61)); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	0 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	118 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_215_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_215_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_215_Update/ca
      -- 
    ca_547_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_215_inst_ack_1, ack => convTranspose_CP_39_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	20 
    -- CP-element group 63: 	24 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_219_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_219_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_219_Sample/rr
      -- 
    rr_555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(63), ack => type_cast_219_inst_req_0); -- 
    convTranspose_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(20) & convTranspose_CP_39_elements(24);
      gj_convTranspose_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_219_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_219_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_219_Sample/ra
      -- 
    ra_556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_219_inst_ack_0, ack => convTranspose_CP_39_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	0 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	118 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_219_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_219_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_219_Update/ca
      -- 
    ca_561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_219_inst_ack_1, ack => convTranspose_CP_39_elements(65)); -- 
    -- CP-element group 66:  join  transition  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	28 
    -- CP-element group 66: 	32 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_256_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_256_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_256_Sample/rr
      -- 
    rr_569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(66), ack => type_cast_256_inst_req_0); -- 
    convTranspose_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(28) & convTranspose_CP_39_elements(32);
      gj_convTranspose_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_256_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_256_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_256_Sample/ra
      -- 
    ra_570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_256_inst_ack_0, ack => convTranspose_CP_39_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	0 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	118 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_256_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_256_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_256_Update/ca
      -- 
    ca_575_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_256_inst_ack_1, ack => convTranspose_CP_39_elements(68)); -- 
    -- CP-element group 69:  join  transition  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	40 
    -- CP-element group 69: 	36 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_260_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_260_Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_260_Sample/rr
      -- 
    rr_583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(69), ack => type_cast_260_inst_req_0); -- 
    convTranspose_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(40) & convTranspose_CP_39_elements(36);
      gj_convTranspose_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_260_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_260_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_260_Sample/ra
      -- 
    ra_584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_260_inst_ack_0, ack => convTranspose_CP_39_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	0 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	118 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_260_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_260_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_260_Update/ca
      -- 
    ca_589_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_260_inst_ack_1, ack => convTranspose_CP_39_elements(71)); -- 
    -- CP-element group 72:  join  transition  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	48 
    -- CP-element group 72: 	44 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_264_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_264_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_264_Sample/rr
      -- 
    rr_597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(72), ack => type_cast_264_inst_req_0); -- 
    convTranspose_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(48) & convTranspose_CP_39_elements(44);
      gj_convTranspose_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_264_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_264_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_264_Sample/ra
      -- 
    ra_598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_264_inst_ack_0, ack => convTranspose_CP_39_elements(73)); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	0 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	118 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_264_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_264_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_264_Update/ca
      -- 
    ca_603_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_264_inst_ack_1, ack => convTranspose_CP_39_elements(74)); -- 
    -- CP-element group 75:  join  transition  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	52 
    -- CP-element group 75: 	56 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_268_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_268_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_268_Sample/rr
      -- 
    rr_611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(75), ack => type_cast_268_inst_req_0); -- 
    convTranspose_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(52) & convTranspose_CP_39_elements(56);
      gj_convTranspose_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_268_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_268_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_268_Sample/ra
      -- 
    ra_612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_268_inst_ack_0, ack => convTranspose_CP_39_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	0 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	118 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_268_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_268_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_268_Update/ca
      -- 
    ca_617_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_268_inst_ack_1, ack => convTranspose_CP_39_elements(77)); -- 
    -- CP-element group 78:  transition  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	54 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (6) 
      -- CP-element group 78: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_286_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_286_update_start_
      -- CP-element group 78: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_286_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_286_Sample/ra
      -- CP-element group 78: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_286_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_286_Update/cr
      -- 
    ra_626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_286_inst_ack_0, ack => convTranspose_CP_39_elements(78)); -- 
    cr_630_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_630_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(78), ack => RPIPE_ConvTranspose_input_pipe_286_inst_req_1); -- 
    -- CP-element group 79:  fork  transition  input  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79: 	82 
    -- CP-element group 79:  members (9) 
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_286_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_286_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_286_Update/ca
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_290_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_290_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_290_Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_299_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_299_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_299_Sample/rr
      -- 
    ca_631_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_286_inst_ack_1, ack => convTranspose_CP_39_elements(79)); -- 
    rr_639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(79), ack => type_cast_290_inst_req_0); -- 
    rr_653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(79), ack => RPIPE_ConvTranspose_input_pipe_299_inst_req_0); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_290_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_290_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_290_Sample/ra
      -- 
    ra_640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_290_inst_ack_0, ack => convTranspose_CP_39_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	0 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	118 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_290_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_290_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_290_Update/ca
      -- 
    ca_645_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_290_inst_ack_1, ack => convTranspose_CP_39_elements(81)); -- 
    -- CP-element group 82:  transition  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	79 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (6) 
      -- CP-element group 82: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_299_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_299_update_start_
      -- CP-element group 82: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_299_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_299_Sample/ra
      -- CP-element group 82: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_299_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_299_Update/cr
      -- 
    ra_654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_299_inst_ack_0, ack => convTranspose_CP_39_elements(82)); -- 
    cr_658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(82), ack => RPIPE_ConvTranspose_input_pipe_299_inst_req_1); -- 
    -- CP-element group 83:  fork  transition  input  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83: 	86 
    -- CP-element group 83:  members (9) 
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_299_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_299_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_299_Update/ca
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_303_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_303_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_303_Sample/rr
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_311_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_311_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_311_Sample/rr
      -- 
    ca_659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_299_inst_ack_1, ack => convTranspose_CP_39_elements(83)); -- 
    rr_667_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_667_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(83), ack => type_cast_303_inst_req_0); -- 
    rr_681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(83), ack => RPIPE_ConvTranspose_input_pipe_311_inst_req_0); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_303_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_303_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_303_Sample/ra
      -- 
    ra_668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_303_inst_ack_0, ack => convTranspose_CP_39_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	0 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	118 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_303_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_303_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_303_Update/ca
      -- 
    ca_673_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_303_inst_ack_1, ack => convTranspose_CP_39_elements(85)); -- 
    -- CP-element group 86:  transition  input  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	83 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (6) 
      -- CP-element group 86: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_311_sample_completed_
      -- CP-element group 86: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_311_update_start_
      -- CP-element group 86: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_311_Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_311_Sample/ra
      -- CP-element group 86: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_311_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_311_Update/cr
      -- 
    ra_682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_311_inst_ack_0, ack => convTranspose_CP_39_elements(86)); -- 
    cr_686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(86), ack => RPIPE_ConvTranspose_input_pipe_311_inst_req_1); -- 
    -- CP-element group 87:  fork  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87: 	90 
    -- CP-element group 87:  members (9) 
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_311_update_completed_
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_311_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_311_Update/ca
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_315_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_315_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_315_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_324_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_324_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_324_Sample/rr
      -- 
    ca_687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_311_inst_ack_1, ack => convTranspose_CP_39_elements(87)); -- 
    rr_695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(87), ack => type_cast_315_inst_req_0); -- 
    rr_709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(87), ack => RPIPE_ConvTranspose_input_pipe_324_inst_req_0); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_315_sample_completed_
      -- CP-element group 88: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_315_Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_315_Sample/ra
      -- 
    ra_696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_315_inst_ack_0, ack => convTranspose_CP_39_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	0 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	118 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_315_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_315_Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_315_Update/ca
      -- 
    ca_701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_315_inst_ack_1, ack => convTranspose_CP_39_elements(89)); -- 
    -- CP-element group 90:  transition  input  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	87 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (6) 
      -- CP-element group 90: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_324_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_324_update_start_
      -- CP-element group 90: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_324_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_324_Sample/ra
      -- CP-element group 90: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_324_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_324_Update/cr
      -- 
    ra_710_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_324_inst_ack_0, ack => convTranspose_CP_39_elements(90)); -- 
    cr_714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(90), ack => RPIPE_ConvTranspose_input_pipe_324_inst_req_1); -- 
    -- CP-element group 91:  fork  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91: 	94 
    -- CP-element group 91:  members (9) 
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_324_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_324_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_324_Update/ca
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_328_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_328_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_328_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_336_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_336_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_336_Sample/rr
      -- 
    ca_715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_324_inst_ack_1, ack => convTranspose_CP_39_elements(91)); -- 
    rr_723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(91), ack => type_cast_328_inst_req_0); -- 
    rr_737_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_737_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(91), ack => RPIPE_ConvTranspose_input_pipe_336_inst_req_0); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_328_sample_completed_
      -- CP-element group 92: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_328_Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_328_Sample/ra
      -- 
    ra_724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_328_inst_ack_0, ack => convTranspose_CP_39_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	0 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	118 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_328_Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_328_update_completed_
      -- CP-element group 93: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_328_Update/ca
      -- 
    ca_729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_328_inst_ack_1, ack => convTranspose_CP_39_elements(93)); -- 
    -- CP-element group 94:  transition  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	91 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (6) 
      -- CP-element group 94: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_336_sample_completed_
      -- CP-element group 94: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_336_update_start_
      -- CP-element group 94: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_336_Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_336_Sample/ra
      -- CP-element group 94: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_336_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_336_Update/cr
      -- 
    ra_738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_336_inst_ack_0, ack => convTranspose_CP_39_elements(94)); -- 
    cr_742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(94), ack => RPIPE_ConvTranspose_input_pipe_336_inst_req_1); -- 
    -- CP-element group 95:  fork  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95: 	98 
    -- CP-element group 95:  members (9) 
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_340_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_340_Sample/rr
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_349_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_349_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_349_Sample/rr
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_336_update_completed_
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_336_Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_336_Update/ca
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_340_sample_start_
      -- 
    ca_743_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_336_inst_ack_1, ack => convTranspose_CP_39_elements(95)); -- 
    rr_751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(95), ack => type_cast_340_inst_req_0); -- 
    rr_765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(95), ack => RPIPE_ConvTranspose_input_pipe_349_inst_req_0); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_340_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_340_Sample/ra
      -- CP-element group 96: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_340_sample_completed_
      -- 
    ra_752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_340_inst_ack_0, ack => convTranspose_CP_39_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	0 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	118 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_340_update_completed_
      -- CP-element group 97: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_340_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_340_Update/ca
      -- 
    ca_757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_340_inst_ack_1, ack => convTranspose_CP_39_elements(97)); -- 
    -- CP-element group 98:  transition  input  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	95 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (6) 
      -- CP-element group 98: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_349_sample_completed_
      -- CP-element group 98: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_349_update_start_
      -- CP-element group 98: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_349_Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_349_Sample/ra
      -- CP-element group 98: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_349_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_349_Update/cr
      -- 
    ra_766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_349_inst_ack_0, ack => convTranspose_CP_39_elements(98)); -- 
    cr_770_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_770_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(98), ack => RPIPE_ConvTranspose_input_pipe_349_inst_req_1); -- 
    -- CP-element group 99:  fork  transition  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: 	102 
    -- CP-element group 99:  members (9) 
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_349_update_completed_
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_349_Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_349_Update/ca
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_353_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_353_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_353_Sample/rr
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_361_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_361_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_361_Sample/rr
      -- 
    ca_771_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_349_inst_ack_1, ack => convTranspose_CP_39_elements(99)); -- 
    rr_779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(99), ack => type_cast_353_inst_req_0); -- 
    rr_793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(99), ack => RPIPE_ConvTranspose_input_pipe_361_inst_req_0); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_353_sample_completed_
      -- CP-element group 100: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_353_Sample/$exit
      -- CP-element group 100: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_353_Sample/ra
      -- 
    ra_780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_353_inst_ack_0, ack => convTranspose_CP_39_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	0 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	118 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_353_update_completed_
      -- CP-element group 101: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_353_Update/$exit
      -- CP-element group 101: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_353_Update/ca
      -- 
    ca_785_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_353_inst_ack_1, ack => convTranspose_CP_39_elements(101)); -- 
    -- CP-element group 102:  transition  input  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	99 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102:  members (6) 
      -- CP-element group 102: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_361_sample_completed_
      -- CP-element group 102: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_361_update_start_
      -- CP-element group 102: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_361_Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_361_Sample/ra
      -- CP-element group 102: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_361_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_361_Update/cr
      -- 
    ra_794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_361_inst_ack_0, ack => convTranspose_CP_39_elements(102)); -- 
    cr_798_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_798_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(102), ack => RPIPE_ConvTranspose_input_pipe_361_inst_req_1); -- 
    -- CP-element group 103:  fork  transition  input  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103: 	106 
    -- CP-element group 103:  members (9) 
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_361_update_completed_
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_361_Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_361_Update/ca
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_365_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_365_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_365_Sample/rr
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_374_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_374_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_374_Sample/rr
      -- 
    ca_799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_361_inst_ack_1, ack => convTranspose_CP_39_elements(103)); -- 
    rr_807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(103), ack => type_cast_365_inst_req_0); -- 
    rr_821_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_821_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(103), ack => RPIPE_ConvTranspose_input_pipe_374_inst_req_0); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_365_sample_completed_
      -- CP-element group 104: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_365_Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_365_Sample/ra
      -- 
    ra_808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_365_inst_ack_0, ack => convTranspose_CP_39_elements(104)); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	0 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	118 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_365_update_completed_
      -- CP-element group 105: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_365_Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_365_Update/ca
      -- 
    ca_813_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_365_inst_ack_1, ack => convTranspose_CP_39_elements(105)); -- 
    -- CP-element group 106:  transition  input  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	103 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (6) 
      -- CP-element group 106: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_374_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_374_update_start_
      -- CP-element group 106: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_374_Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_374_Sample/ra
      -- CP-element group 106: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_374_Update/$entry
      -- CP-element group 106: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_374_Update/cr
      -- 
    ra_822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_374_inst_ack_0, ack => convTranspose_CP_39_elements(106)); -- 
    cr_826_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_826_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(106), ack => RPIPE_ConvTranspose_input_pipe_374_inst_req_1); -- 
    -- CP-element group 107:  fork  transition  input  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107: 	110 
    -- CP-element group 107:  members (9) 
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_374_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_374_Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_374_Update/ca
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_378_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_378_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_378_Sample/rr
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_386_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_386_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_386_Sample/rr
      -- 
    ca_827_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_374_inst_ack_1, ack => convTranspose_CP_39_elements(107)); -- 
    rr_835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(107), ack => type_cast_378_inst_req_0); -- 
    rr_849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(107), ack => RPIPE_ConvTranspose_input_pipe_386_inst_req_0); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_378_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_378_Sample/$exit
      -- CP-element group 108: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_378_Sample/ra
      -- 
    ra_836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_378_inst_ack_0, ack => convTranspose_CP_39_elements(108)); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	0 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	118 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_378_update_completed_
      -- CP-element group 109: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_378_Update/$exit
      -- CP-element group 109: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_378_Update/ca
      -- 
    ca_841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_378_inst_ack_1, ack => convTranspose_CP_39_elements(109)); -- 
    -- CP-element group 110:  transition  input  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	107 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (6) 
      -- CP-element group 110: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_386_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_386_update_start_
      -- CP-element group 110: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_386_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_386_Sample/ra
      -- CP-element group 110: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_386_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_386_Update/cr
      -- 
    ra_850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_386_inst_ack_0, ack => convTranspose_CP_39_elements(110)); -- 
    cr_854_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_854_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(110), ack => RPIPE_ConvTranspose_input_pipe_386_inst_req_1); -- 
    -- CP-element group 111:  fork  transition  input  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111: 	114 
    -- CP-element group 111:  members (9) 
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_386_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_386_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_386_Update/ca
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_390_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_390_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_390_Sample/rr
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_399_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_399_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_399_Sample/rr
      -- 
    ca_855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_386_inst_ack_1, ack => convTranspose_CP_39_elements(111)); -- 
    rr_863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(111), ack => type_cast_390_inst_req_0); -- 
    rr_877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(111), ack => RPIPE_ConvTranspose_input_pipe_399_inst_req_0); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_390_sample_completed_
      -- CP-element group 112: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_390_Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_390_Sample/ra
      -- 
    ra_864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_390_inst_ack_0, ack => convTranspose_CP_39_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	0 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	118 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_390_update_completed_
      -- CP-element group 113: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_390_Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_390_Update/ca
      -- 
    ca_869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_390_inst_ack_1, ack => convTranspose_CP_39_elements(113)); -- 
    -- CP-element group 114:  transition  input  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	111 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (6) 
      -- CP-element group 114: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_399_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_399_update_start_
      -- CP-element group 114: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_399_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_399_Sample/ra
      -- CP-element group 114: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_399_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_399_Update/cr
      -- 
    ra_878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_399_inst_ack_0, ack => convTranspose_CP_39_elements(114)); -- 
    cr_882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(114), ack => RPIPE_ConvTranspose_input_pipe_399_inst_req_1); -- 
    -- CP-element group 115:  transition  input  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (6) 
      -- CP-element group 115: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_399_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_399_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_399_Update/ca
      -- CP-element group 115: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_403_sample_start_
      -- CP-element group 115: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_403_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_403_Sample/rr
      -- 
    ca_883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_399_inst_ack_1, ack => convTranspose_CP_39_elements(115)); -- 
    rr_891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(115), ack => type_cast_403_inst_req_0); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_403_sample_completed_
      -- CP-element group 116: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_403_Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_403_Sample/ra
      -- 
    ra_892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_403_inst_ack_0, ack => convTranspose_CP_39_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	0 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_403_update_completed_
      -- CP-element group 117: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_403_Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_403_Update/ca
      -- 
    ca_897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_403_inst_ack_1, ack => convTranspose_CP_39_elements(117)); -- 
    -- CP-element group 118:  branch  join  transition  place  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	59 
    -- CP-element group 118: 	62 
    -- CP-element group 118: 	65 
    -- CP-element group 118: 	68 
    -- CP-element group 118: 	71 
    -- CP-element group 118: 	74 
    -- CP-element group 118: 	77 
    -- CP-element group 118: 	81 
    -- CP-element group 118: 	85 
    -- CP-element group 118: 	89 
    -- CP-element group 118: 	93 
    -- CP-element group 118: 	97 
    -- CP-element group 118: 	101 
    -- CP-element group 118: 	105 
    -- CP-element group 118: 	109 
    -- CP-element group 118: 	113 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118: 	120 
    -- CP-element group 118:  members (10) 
      -- CP-element group 118: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416__exit__
      -- CP-element group 118: 	 branch_block_stmt_33/if_stmt_417__entry__
      -- CP-element group 118: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/$exit
      -- CP-element group 118: 	 branch_block_stmt_33/if_stmt_417_dead_link/$entry
      -- CP-element group 118: 	 branch_block_stmt_33/if_stmt_417_eval_test/$entry
      -- CP-element group 118: 	 branch_block_stmt_33/if_stmt_417_eval_test/$exit
      -- CP-element group 118: 	 branch_block_stmt_33/if_stmt_417_eval_test/branch_req
      -- CP-element group 118: 	 branch_block_stmt_33/R_cmp514_418_place
      -- CP-element group 118: 	 branch_block_stmt_33/if_stmt_417_if_link/$entry
      -- CP-element group 118: 	 branch_block_stmt_33/if_stmt_417_else_link/$entry
      -- 
    branch_req_905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(118), ack => if_stmt_417_branch_req_0); -- 
    convTranspose_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(59) & convTranspose_CP_39_elements(62) & convTranspose_CP_39_elements(65) & convTranspose_CP_39_elements(68) & convTranspose_CP_39_elements(71) & convTranspose_CP_39_elements(74) & convTranspose_CP_39_elements(77) & convTranspose_CP_39_elements(81) & convTranspose_CP_39_elements(85) & convTranspose_CP_39_elements(89) & convTranspose_CP_39_elements(93) & convTranspose_CP_39_elements(97) & convTranspose_CP_39_elements(101) & convTranspose_CP_39_elements(105) & convTranspose_CP_39_elements(109) & convTranspose_CP_39_elements(113) & convTranspose_CP_39_elements(117);
      gj_convTranspose_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	123 
    -- CP-element group 119: 	124 
    -- CP-element group 119:  members (18) 
      -- CP-element group 119: 	 branch_block_stmt_33/merge_stmt_438__exit__
      -- CP-element group 119: 	 branch_block_stmt_33/assign_stmt_444_to_assign_stmt_467__entry__
      -- CP-element group 119: 	 branch_block_stmt_33/if_stmt_417_if_link/$exit
      -- CP-element group 119: 	 branch_block_stmt_33/if_stmt_417_if_link/if_choice_transition
      -- CP-element group 119: 	 branch_block_stmt_33/entry_bbx_xnph516
      -- CP-element group 119: 	 branch_block_stmt_33/assign_stmt_444_to_assign_stmt_467/$entry
      -- CP-element group 119: 	 branch_block_stmt_33/assign_stmt_444_to_assign_stmt_467/type_cast_453_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_33/assign_stmt_444_to_assign_stmt_467/type_cast_453_update_start_
      -- CP-element group 119: 	 branch_block_stmt_33/assign_stmt_444_to_assign_stmt_467/type_cast_453_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_33/assign_stmt_444_to_assign_stmt_467/type_cast_453_Sample/rr
      -- CP-element group 119: 	 branch_block_stmt_33/assign_stmt_444_to_assign_stmt_467/type_cast_453_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_33/assign_stmt_444_to_assign_stmt_467/type_cast_453_Update/cr
      -- CP-element group 119: 	 branch_block_stmt_33/entry_bbx_xnph516_PhiReq/$entry
      -- CP-element group 119: 	 branch_block_stmt_33/entry_bbx_xnph516_PhiReq/$exit
      -- CP-element group 119: 	 branch_block_stmt_33/merge_stmt_438_PhiReqMerge
      -- CP-element group 119: 	 branch_block_stmt_33/merge_stmt_438_PhiAck/$entry
      -- CP-element group 119: 	 branch_block_stmt_33/merge_stmt_438_PhiAck/$exit
      -- CP-element group 119: 	 branch_block_stmt_33/merge_stmt_438_PhiAck/dummy
      -- 
    if_choice_transition_910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_417_branch_ack_1, ack => convTranspose_CP_39_elements(119)); -- 
    rr_949_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_949_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(119), ack => type_cast_453_inst_req_0); -- 
    cr_954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(119), ack => type_cast_453_inst_req_1); -- 
    -- CP-element group 120:  transition  place  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	118 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	472 
    -- CP-element group 120:  members (5) 
      -- CP-element group 120: 	 branch_block_stmt_33/if_stmt_417_else_link/$exit
      -- CP-element group 120: 	 branch_block_stmt_33/if_stmt_417_else_link/else_choice_transition
      -- CP-element group 120: 	 branch_block_stmt_33/entry_forx_xcond190x_xpreheader
      -- CP-element group 120: 	 branch_block_stmt_33/entry_forx_xcond190x_xpreheader_PhiReq/$entry
      -- CP-element group 120: 	 branch_block_stmt_33/entry_forx_xcond190x_xpreheader_PhiReq/$exit
      -- 
    else_choice_transition_914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_417_branch_ack_0, ack => convTranspose_CP_39_elements(120)); -- 
    -- CP-element group 121:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	472 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	167 
    -- CP-element group 121: 	168 
    -- CP-element group 121:  members (18) 
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_645_to_assign_stmt_674/type_cast_660_update_start_
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_645_to_assign_stmt_674/type_cast_660_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_33/merge_stmt_639__exit__
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_645_to_assign_stmt_674__entry__
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_645_to_assign_stmt_674/type_cast_660_Update/$entry
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_645_to_assign_stmt_674/$entry
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_645_to_assign_stmt_674/type_cast_660_Sample/rr
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_645_to_assign_stmt_674/type_cast_660_Sample/$entry
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_645_to_assign_stmt_674/type_cast_660_Update/cr
      -- CP-element group 121: 	 branch_block_stmt_33/if_stmt_432_if_link/$exit
      -- CP-element group 121: 	 branch_block_stmt_33/if_stmt_432_if_link/if_choice_transition
      -- CP-element group 121: 	 branch_block_stmt_33/forx_xcond190x_xpreheader_bbx_xnph512
      -- CP-element group 121: 	 branch_block_stmt_33/forx_xcond190x_xpreheader_bbx_xnph512_PhiReq/$entry
      -- CP-element group 121: 	 branch_block_stmt_33/forx_xcond190x_xpreheader_bbx_xnph512_PhiReq/$exit
      -- CP-element group 121: 	 branch_block_stmt_33/merge_stmt_639_PhiReqMerge
      -- CP-element group 121: 	 branch_block_stmt_33/merge_stmt_639_PhiAck/$entry
      -- CP-element group 121: 	 branch_block_stmt_33/merge_stmt_639_PhiAck/$exit
      -- CP-element group 121: 	 branch_block_stmt_33/merge_stmt_639_PhiAck/dummy
      -- 
    if_choice_transition_932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_432_branch_ack_1, ack => convTranspose_CP_39_elements(121)); -- 
    rr_1308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(121), ack => type_cast_660_inst_req_0); -- 
    cr_1313_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1313_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(121), ack => type_cast_660_inst_req_1); -- 
    -- CP-element group 122:  transition  place  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	472 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	485 
    -- CP-element group 122:  members (5) 
      -- CP-element group 122: 	 branch_block_stmt_33/if_stmt_432_else_link/$exit
      -- CP-element group 122: 	 branch_block_stmt_33/if_stmt_432_else_link/else_choice_transition
      -- CP-element group 122: 	 branch_block_stmt_33/forx_xcond190x_xpreheader_forx_xend250
      -- CP-element group 122: 	 branch_block_stmt_33/forx_xcond190x_xpreheader_forx_xend250_PhiReq/$entry
      -- CP-element group 122: 	 branch_block_stmt_33/forx_xcond190x_xpreheader_forx_xend250_PhiReq/$exit
      -- 
    else_choice_transition_936_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_432_branch_ack_0, ack => convTranspose_CP_39_elements(122)); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	119 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_33/assign_stmt_444_to_assign_stmt_467/type_cast_453_sample_completed_
      -- CP-element group 123: 	 branch_block_stmt_33/assign_stmt_444_to_assign_stmt_467/type_cast_453_Sample/$exit
      -- CP-element group 123: 	 branch_block_stmt_33/assign_stmt_444_to_assign_stmt_467/type_cast_453_Sample/ra
      -- 
    ra_950_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_453_inst_ack_0, ack => convTranspose_CP_39_elements(123)); -- 
    -- CP-element group 124:  transition  place  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	119 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	473 
    -- CP-element group 124:  members (9) 
      -- CP-element group 124: 	 branch_block_stmt_33/assign_stmt_444_to_assign_stmt_467__exit__
      -- CP-element group 124: 	 branch_block_stmt_33/bbx_xnph516_forx_xbody
      -- CP-element group 124: 	 branch_block_stmt_33/assign_stmt_444_to_assign_stmt_467/$exit
      -- CP-element group 124: 	 branch_block_stmt_33/assign_stmt_444_to_assign_stmt_467/type_cast_453_update_completed_
      -- CP-element group 124: 	 branch_block_stmt_33/assign_stmt_444_to_assign_stmt_467/type_cast_453_Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_33/assign_stmt_444_to_assign_stmt_467/type_cast_453_Update/ca
      -- CP-element group 124: 	 branch_block_stmt_33/bbx_xnph516_forx_xbody_PhiReq/$entry
      -- CP-element group 124: 	 branch_block_stmt_33/bbx_xnph516_forx_xbody_PhiReq/phi_stmt_470/$entry
      -- CP-element group 124: 	 branch_block_stmt_33/bbx_xnph516_forx_xbody_PhiReq/phi_stmt_470/phi_stmt_470_sources/$entry
      -- 
    ca_955_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_453_inst_ack_1, ack => convTranspose_CP_39_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	478 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	164 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_final_index_sum_regn_sample_complete
      -- CP-element group 125: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_final_index_sum_regn_Sample/$exit
      -- CP-element group 125: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_final_index_sum_regn_Sample/ack
      -- 
    ack_984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_482_index_offset_ack_0, ack => convTranspose_CP_39_elements(125)); -- 
    -- CP-element group 126:  transition  input  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	478 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (11) 
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/addr_of_483_sample_start_
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_root_address_calculated
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_offset_calculated
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_final_index_sum_regn_Update/$exit
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_final_index_sum_regn_Update/ack
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_base_plus_offset/$entry
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_base_plus_offset/$exit
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_base_plus_offset/sum_rename_req
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_base_plus_offset/sum_rename_ack
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/addr_of_483_request/$entry
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/addr_of_483_request/req
      -- 
    ack_989_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_482_index_offset_ack_1, ack => convTranspose_CP_39_elements(126)); -- 
    req_998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(126), ack => addr_of_483_final_reg_req_0); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/addr_of_483_sample_completed_
      -- CP-element group 127: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/addr_of_483_request/$exit
      -- CP-element group 127: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/addr_of_483_request/ack
      -- 
    ack_999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_483_final_reg_ack_0, ack => convTranspose_CP_39_elements(127)); -- 
    -- CP-element group 128:  fork  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	478 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	161 
    -- CP-element group 128:  members (19) 
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_base_plus_offset/sum_rename_req
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_word_addrgen/root_register_ack
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_word_addrgen/root_register_req
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_word_addrgen/$exit
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_word_addrgen/$entry
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_base_plus_offset/sum_rename_ack
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_base_plus_offset/$exit
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_base_plus_offset/$entry
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_base_addr_resize/base_resize_ack
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_base_addr_resize/base_resize_req
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_base_addr_resize/$exit
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_base_addr_resize/$entry
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_base_address_resized
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_root_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_word_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_base_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/addr_of_483_update_completed_
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/addr_of_483_complete/$exit
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/addr_of_483_complete/ack
      -- 
    ack_1004_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_483_final_reg_ack_1, ack => convTranspose_CP_39_elements(128)); -- 
    -- CP-element group 129:  transition  input  output  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	478 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (6) 
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_486_sample_completed_
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_486_update_start_
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_486_Sample/$exit
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_486_Sample/ra
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_486_Update/$entry
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_486_Update/cr
      -- 
    ra_1013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_486_inst_ack_0, ack => convTranspose_CP_39_elements(129)); -- 
    cr_1017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(129), ack => RPIPE_ConvTranspose_input_pipe_486_inst_req_1); -- 
    -- CP-element group 130:  fork  transition  input  output  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130: 	133 
    -- CP-element group 130:  members (9) 
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_486_update_completed_
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_486_Update/$exit
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_486_Update/ca
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_490_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_490_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_490_Sample/rr
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_499_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_499_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_499_Sample/rr
      -- 
    ca_1018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_486_inst_ack_1, ack => convTranspose_CP_39_elements(130)); -- 
    rr_1026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(130), ack => type_cast_490_inst_req_0); -- 
    rr_1040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(130), ack => RPIPE_ConvTranspose_input_pipe_499_inst_req_0); -- 
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_490_sample_completed_
      -- CP-element group 131: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_490_Sample/$exit
      -- CP-element group 131: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_490_Sample/ra
      -- 
    ra_1027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_490_inst_ack_0, ack => convTranspose_CP_39_elements(131)); -- 
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	478 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	161 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_490_update_completed_
      -- CP-element group 132: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_490_Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_490_Update/ca
      -- 
    ca_1032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_490_inst_ack_1, ack => convTranspose_CP_39_elements(132)); -- 
    -- CP-element group 133:  transition  input  output  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	130 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133:  members (6) 
      -- CP-element group 133: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_499_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_499_update_start_
      -- CP-element group 133: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_499_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_499_Sample/ra
      -- CP-element group 133: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_499_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_499_Update/cr
      -- 
    ra_1041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_499_inst_ack_0, ack => convTranspose_CP_39_elements(133)); -- 
    cr_1045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(133), ack => RPIPE_ConvTranspose_input_pipe_499_inst_req_1); -- 
    -- CP-element group 134:  fork  transition  input  output  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134: 	137 
    -- CP-element group 134:  members (9) 
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_499_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_499_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_499_Update/ca
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_503_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_503_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_503_Sample/rr
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_517_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_517_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_517_Sample/rr
      -- 
    ca_1046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_499_inst_ack_1, ack => convTranspose_CP_39_elements(134)); -- 
    rr_1054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(134), ack => type_cast_503_inst_req_0); -- 
    rr_1068_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1068_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(134), ack => RPIPE_ConvTranspose_input_pipe_517_inst_req_0); -- 
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	134 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_503_sample_completed_
      -- CP-element group 135: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_503_Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_503_Sample/ra
      -- 
    ra_1055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_503_inst_ack_0, ack => convTranspose_CP_39_elements(135)); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	478 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	161 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_503_update_completed_
      -- CP-element group 136: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_503_Update/$exit
      -- CP-element group 136: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_503_Update/ca
      -- 
    ca_1060_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_503_inst_ack_1, ack => convTranspose_CP_39_elements(136)); -- 
    -- CP-element group 137:  transition  input  output  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	134 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137:  members (6) 
      -- CP-element group 137: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_517_sample_completed_
      -- CP-element group 137: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_517_update_start_
      -- CP-element group 137: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_517_Sample/$exit
      -- CP-element group 137: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_517_Sample/ra
      -- CP-element group 137: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_517_Update/$entry
      -- CP-element group 137: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_517_Update/cr
      -- 
    ra_1069_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_517_inst_ack_0, ack => convTranspose_CP_39_elements(137)); -- 
    cr_1073_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1073_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(137), ack => RPIPE_ConvTranspose_input_pipe_517_inst_req_1); -- 
    -- CP-element group 138:  fork  transition  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	139 
    -- CP-element group 138: 	141 
    -- CP-element group 138:  members (9) 
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_535_Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_535_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_521_Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_535_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_517_update_completed_
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_517_Update/$exit
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_517_Update/ca
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_521_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_521_Sample/$entry
      -- 
    ca_1074_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_517_inst_ack_1, ack => convTranspose_CP_39_elements(138)); -- 
    rr_1082_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1082_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(138), ack => type_cast_521_inst_req_0); -- 
    rr_1096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(138), ack => RPIPE_ConvTranspose_input_pipe_535_inst_req_0); -- 
    -- CP-element group 139:  transition  input  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	138 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_521_Sample/ra
      -- CP-element group 139: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_521_Sample/$exit
      -- CP-element group 139: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_521_sample_completed_
      -- 
    ra_1083_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_521_inst_ack_0, ack => convTranspose_CP_39_elements(139)); -- 
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	478 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	161 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_521_Update/ca
      -- CP-element group 140: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_521_Update/$exit
      -- CP-element group 140: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_521_update_completed_
      -- 
    ca_1088_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_521_inst_ack_1, ack => convTranspose_CP_39_elements(140)); -- 
    -- CP-element group 141:  transition  input  output  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	138 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	142 
    -- CP-element group 141:  members (6) 
      -- CP-element group 141: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_535_Update/cr
      -- CP-element group 141: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_535_Update/$entry
      -- CP-element group 141: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_535_Sample/ra
      -- CP-element group 141: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_535_Sample/$exit
      -- CP-element group 141: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_535_update_start_
      -- CP-element group 141: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_535_sample_completed_
      -- 
    ra_1097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_535_inst_ack_0, ack => convTranspose_CP_39_elements(141)); -- 
    cr_1101_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1101_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(141), ack => RPIPE_ConvTranspose_input_pipe_535_inst_req_1); -- 
    -- CP-element group 142:  fork  transition  input  output  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	141 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	143 
    -- CP-element group 142: 	145 
    -- CP-element group 142:  members (9) 
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_539_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_535_Update/ca
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_535_Update/$exit
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_535_update_completed_
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_553_Sample/rr
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_553_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_553_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_539_Sample/rr
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_539_Sample/$entry
      -- 
    ca_1102_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_535_inst_ack_1, ack => convTranspose_CP_39_elements(142)); -- 
    rr_1110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(142), ack => type_cast_539_inst_req_0); -- 
    rr_1124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(142), ack => RPIPE_ConvTranspose_input_pipe_553_inst_req_0); -- 
    -- CP-element group 143:  transition  input  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	142 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_539_sample_completed_
      -- CP-element group 143: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_539_Sample/ra
      -- CP-element group 143: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_539_Sample/$exit
      -- 
    ra_1111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_539_inst_ack_0, ack => convTranspose_CP_39_elements(143)); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	478 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	161 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_539_update_completed_
      -- CP-element group 144: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_539_Update/ca
      -- CP-element group 144: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_539_Update/$exit
      -- 
    ca_1116_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_539_inst_ack_1, ack => convTranspose_CP_39_elements(144)); -- 
    -- CP-element group 145:  transition  input  output  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	142 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145:  members (6) 
      -- CP-element group 145: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_553_Update/cr
      -- CP-element group 145: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_553_Update/$entry
      -- CP-element group 145: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_553_Sample/ra
      -- CP-element group 145: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_553_Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_553_update_start_
      -- CP-element group 145: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_553_sample_completed_
      -- 
    ra_1125_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_553_inst_ack_0, ack => convTranspose_CP_39_elements(145)); -- 
    cr_1129_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1129_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(145), ack => RPIPE_ConvTranspose_input_pipe_553_inst_req_1); -- 
    -- CP-element group 146:  fork  transition  input  output  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	145 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	147 
    -- CP-element group 146: 	149 
    -- CP-element group 146:  members (9) 
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_571_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_571_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_571_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_557_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_557_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_557_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_553_Update/ca
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_553_Update/$exit
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_553_update_completed_
      -- 
    ca_1130_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_553_inst_ack_1, ack => convTranspose_CP_39_elements(146)); -- 
    rr_1138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(146), ack => type_cast_557_inst_req_0); -- 
    rr_1152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(146), ack => RPIPE_ConvTranspose_input_pipe_571_inst_req_0); -- 
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	146 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_557_Sample/ra
      -- CP-element group 147: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_557_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_557_sample_completed_
      -- 
    ra_1139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_557_inst_ack_0, ack => convTranspose_CP_39_elements(147)); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	478 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	161 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_557_Update/ca
      -- CP-element group 148: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_557_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_557_update_completed_
      -- 
    ca_1144_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_557_inst_ack_1, ack => convTranspose_CP_39_elements(148)); -- 
    -- CP-element group 149:  transition  input  output  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	146 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	150 
    -- CP-element group 149:  members (6) 
      -- CP-element group 149: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_571_Sample/ra
      -- CP-element group 149: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_571_Update/cr
      -- CP-element group 149: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_571_Update/$entry
      -- CP-element group 149: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_571_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_571_update_start_
      -- CP-element group 149: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_571_sample_completed_
      -- 
    ra_1153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_571_inst_ack_0, ack => convTranspose_CP_39_elements(149)); -- 
    cr_1157_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1157_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(149), ack => RPIPE_ConvTranspose_input_pipe_571_inst_req_1); -- 
    -- CP-element group 150:  fork  transition  input  output  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	149 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	151 
    -- CP-element group 150: 	153 
    -- CP-element group 150:  members (9) 
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_589_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_589_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_589_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_575_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_575_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_575_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_571_Update/ca
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_571_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_571_update_completed_
      -- 
    ca_1158_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_571_inst_ack_1, ack => convTranspose_CP_39_elements(150)); -- 
    rr_1166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(150), ack => type_cast_575_inst_req_0); -- 
    rr_1180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(150), ack => RPIPE_ConvTranspose_input_pipe_589_inst_req_0); -- 
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	150 
    -- CP-element group 151: successors 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_575_Sample/ra
      -- CP-element group 151: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_575_sample_completed_
      -- CP-element group 151: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_575_Sample/$exit
      -- 
    ra_1167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_575_inst_ack_0, ack => convTranspose_CP_39_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	478 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	161 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_575_Update/ca
      -- CP-element group 152: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_575_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_575_update_completed_
      -- 
    ca_1172_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_575_inst_ack_1, ack => convTranspose_CP_39_elements(152)); -- 
    -- CP-element group 153:  transition  input  output  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	150 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153:  members (6) 
      -- CP-element group 153: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_589_Update/cr
      -- CP-element group 153: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_589_Update/$entry
      -- CP-element group 153: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_589_Sample/ra
      -- CP-element group 153: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_589_Sample/$exit
      -- CP-element group 153: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_589_update_start_
      -- CP-element group 153: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_589_sample_completed_
      -- 
    ra_1181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_589_inst_ack_0, ack => convTranspose_CP_39_elements(153)); -- 
    cr_1185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(153), ack => RPIPE_ConvTranspose_input_pipe_589_inst_req_1); -- 
    -- CP-element group 154:  fork  transition  input  output  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154: 	157 
    -- CP-element group 154:  members (9) 
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_589_Update/ca
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_589_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_589_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_607_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_607_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_607_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_593_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_593_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_593_sample_start_
      -- 
    ca_1186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_589_inst_ack_1, ack => convTranspose_CP_39_elements(154)); -- 
    rr_1208_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1208_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(154), ack => RPIPE_ConvTranspose_input_pipe_607_inst_req_0); -- 
    rr_1194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(154), ack => type_cast_593_inst_req_0); -- 
    -- CP-element group 155:  transition  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_593_Sample/ra
      -- CP-element group 155: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_593_Sample/$exit
      -- CP-element group 155: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_593_sample_completed_
      -- 
    ra_1195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_593_inst_ack_0, ack => convTranspose_CP_39_elements(155)); -- 
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	478 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	161 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_593_Update/ca
      -- CP-element group 156: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_593_Update/$exit
      -- CP-element group 156: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_593_update_completed_
      -- 
    ca_1200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_593_inst_ack_1, ack => convTranspose_CP_39_elements(156)); -- 
    -- CP-element group 157:  transition  input  output  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	154 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	158 
    -- CP-element group 157:  members (6) 
      -- CP-element group 157: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_607_Update/cr
      -- CP-element group 157: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_607_Update/$entry
      -- CP-element group 157: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_607_Sample/ra
      -- CP-element group 157: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_607_Sample/$exit
      -- CP-element group 157: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_607_update_start_
      -- CP-element group 157: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_607_sample_completed_
      -- 
    ra_1209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_607_inst_ack_0, ack => convTranspose_CP_39_elements(157)); -- 
    cr_1213_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1213_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(157), ack => RPIPE_ConvTranspose_input_pipe_607_inst_req_1); -- 
    -- CP-element group 158:  transition  input  output  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	157 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	159 
    -- CP-element group 158:  members (6) 
      -- CP-element group 158: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_611_sample_start_
      -- CP-element group 158: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_607_Update/ca
      -- CP-element group 158: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_607_Update/$exit
      -- CP-element group 158: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_607_update_completed_
      -- CP-element group 158: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_611_Sample/rr
      -- CP-element group 158: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_611_Sample/$entry
      -- 
    ca_1214_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_607_inst_ack_1, ack => convTranspose_CP_39_elements(158)); -- 
    rr_1222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(158), ack => type_cast_611_inst_req_0); -- 
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	158 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_611_sample_completed_
      -- CP-element group 159: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_611_Sample/ra
      -- CP-element group 159: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_611_Sample/$exit
      -- 
    ra_1223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_611_inst_ack_0, ack => convTranspose_CP_39_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	478 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	161 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_611_update_completed_
      -- CP-element group 160: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_611_Update/ca
      -- CP-element group 160: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_611_Update/$exit
      -- 
    ca_1228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_611_inst_ack_1, ack => convTranspose_CP_39_elements(160)); -- 
    -- CP-element group 161:  join  transition  output  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	156 
    -- CP-element group 161: 	160 
    -- CP-element group 161: 	128 
    -- CP-element group 161: 	132 
    -- CP-element group 161: 	136 
    -- CP-element group 161: 	140 
    -- CP-element group 161: 	144 
    -- CP-element group 161: 	148 
    -- CP-element group 161: 	152 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161:  members (9) 
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_Sample/word_access_start/word_0/$entry
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_Sample/word_access_start/$entry
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_Sample/ptr_deref_619_Split/split_ack
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_Sample/ptr_deref_619_Split/split_req
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_Sample/ptr_deref_619_Split/$exit
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_Sample/ptr_deref_619_Split/$entry
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_Sample/$entry
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_sample_start_
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_Sample/word_access_start/word_0/rr
      -- 
    rr_1266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(161), ack => ptr_deref_619_store_0_req_0); -- 
    convTranspose_cp_element_group_161: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_161"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(156) & convTranspose_CP_39_elements(160) & convTranspose_CP_39_elements(128) & convTranspose_CP_39_elements(132) & convTranspose_CP_39_elements(136) & convTranspose_CP_39_elements(140) & convTranspose_CP_39_elements(144) & convTranspose_CP_39_elements(148) & convTranspose_CP_39_elements(152);
      gj_convTranspose_cp_element_group_161 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(161), clk => clk, reset => reset); --
    end block;
    -- CP-element group 162:  transition  input  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	161 
    -- CP-element group 162: successors 
    -- CP-element group 162:  members (5) 
      -- CP-element group 162: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_Sample/word_access_start/word_0/$exit
      -- CP-element group 162: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_Sample/word_access_start/$exit
      -- CP-element group 162: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_Sample/$exit
      -- CP-element group 162: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_sample_completed_
      -- CP-element group 162: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_Sample/word_access_start/word_0/ra
      -- 
    ra_1267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_619_store_0_ack_0, ack => convTranspose_CP_39_elements(162)); -- 
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	478 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	164 
    -- CP-element group 163:  members (5) 
      -- CP-element group 163: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_Update/word_access_complete/word_0/ca
      -- CP-element group 163: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_update_completed_
      -- CP-element group 163: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_Update/word_access_complete/word_0/$exit
      -- CP-element group 163: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_Update/word_access_complete/$exit
      -- CP-element group 163: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_Update/$exit
      -- 
    ca_1278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_619_store_0_ack_1, ack => convTranspose_CP_39_elements(163)); -- 
    -- CP-element group 164:  branch  join  transition  place  output  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	163 
    -- CP-element group 164: 	125 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	165 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (10) 
      -- CP-element group 164: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632__exit__
      -- CP-element group 164: 	 branch_block_stmt_33/if_stmt_633__entry__
      -- CP-element group 164: 	 branch_block_stmt_33/if_stmt_633_else_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_33/if_stmt_633_if_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_33/R_exitcond3_634_place
      -- CP-element group 164: 	 branch_block_stmt_33/if_stmt_633_eval_test/branch_req
      -- CP-element group 164: 	 branch_block_stmt_33/if_stmt_633_eval_test/$exit
      -- CP-element group 164: 	 branch_block_stmt_33/if_stmt_633_eval_test/$entry
      -- CP-element group 164: 	 branch_block_stmt_33/if_stmt_633_dead_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/$exit
      -- 
    branch_req_1286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(164), ack => if_stmt_633_branch_req_0); -- 
    convTranspose_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(163) & convTranspose_CP_39_elements(125);
      gj_convTranspose_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  merge  transition  place  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	164 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	472 
    -- CP-element group 165:  members (13) 
      -- CP-element group 165: 	 branch_block_stmt_33/merge_stmt_423__exit__
      -- CP-element group 165: 	 branch_block_stmt_33/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader
      -- CP-element group 165: 	 branch_block_stmt_33/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit
      -- CP-element group 165: 	 branch_block_stmt_33/if_stmt_633_if_link/if_choice_transition
      -- CP-element group 165: 	 branch_block_stmt_33/if_stmt_633_if_link/$exit
      -- CP-element group 165: 	 branch_block_stmt_33/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit_PhiReq/$entry
      -- CP-element group 165: 	 branch_block_stmt_33/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit_PhiReq/$exit
      -- CP-element group 165: 	 branch_block_stmt_33/merge_stmt_423_PhiReqMerge
      -- CP-element group 165: 	 branch_block_stmt_33/merge_stmt_423_PhiAck/$entry
      -- CP-element group 165: 	 branch_block_stmt_33/merge_stmt_423_PhiAck/$exit
      -- CP-element group 165: 	 branch_block_stmt_33/merge_stmt_423_PhiAck/dummy
      -- CP-element group 165: 	 branch_block_stmt_33/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader_PhiReq/$entry
      -- CP-element group 165: 	 branch_block_stmt_33/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader_PhiReq/$exit
      -- 
    if_choice_transition_1291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_633_branch_ack_1, ack => convTranspose_CP_39_elements(165)); -- 
    -- CP-element group 166:  fork  transition  place  input  output  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	474 
    -- CP-element group 166: 	475 
    -- CP-element group 166:  members (12) 
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody_forx_xbody
      -- CP-element group 166: 	 branch_block_stmt_33/if_stmt_633_else_link/else_choice_transition
      -- CP-element group 166: 	 branch_block_stmt_33/if_stmt_633_else_link/$exit
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_470/$entry
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_470/phi_stmt_470_sources/$entry
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_470/phi_stmt_470_sources/type_cast_476/$entry
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_470/phi_stmt_470_sources/type_cast_476/SplitProtocol/$entry
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_470/phi_stmt_470_sources/type_cast_476/SplitProtocol/Sample/$entry
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_470/phi_stmt_470_sources/type_cast_476/SplitProtocol/Sample/rr
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_470/phi_stmt_470_sources/type_cast_476/SplitProtocol/Update/$entry
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_470/phi_stmt_470_sources/type_cast_476/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1295_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_633_branch_ack_0, ack => convTranspose_CP_39_elements(166)); -- 
    rr_3525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(166), ack => type_cast_476_inst_req_0); -- 
    cr_3530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(166), ack => type_cast_476_inst_req_1); -- 
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	121 
    -- CP-element group 167: successors 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_33/assign_stmt_645_to_assign_stmt_674/type_cast_660_sample_completed_
      -- CP-element group 167: 	 branch_block_stmt_33/assign_stmt_645_to_assign_stmt_674/type_cast_660_Sample/ra
      -- CP-element group 167: 	 branch_block_stmt_33/assign_stmt_645_to_assign_stmt_674/type_cast_660_Sample/$exit
      -- 
    ra_1309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_660_inst_ack_0, ack => convTranspose_CP_39_elements(167)); -- 
    -- CP-element group 168:  transition  place  input  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	121 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	479 
    -- CP-element group 168:  members (9) 
      -- CP-element group 168: 	 branch_block_stmt_33/assign_stmt_645_to_assign_stmt_674/type_cast_660_Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_33/assign_stmt_645_to_assign_stmt_674__exit__
      -- CP-element group 168: 	 branch_block_stmt_33/bbx_xnph512_forx_xbody196
      -- CP-element group 168: 	 branch_block_stmt_33/assign_stmt_645_to_assign_stmt_674/$exit
      -- CP-element group 168: 	 branch_block_stmt_33/assign_stmt_645_to_assign_stmt_674/type_cast_660_update_completed_
      -- CP-element group 168: 	 branch_block_stmt_33/assign_stmt_645_to_assign_stmt_674/type_cast_660_Update/ca
      -- CP-element group 168: 	 branch_block_stmt_33/bbx_xnph512_forx_xbody196_PhiReq/$entry
      -- CP-element group 168: 	 branch_block_stmt_33/bbx_xnph512_forx_xbody196_PhiReq/phi_stmt_677/$entry
      -- CP-element group 168: 	 branch_block_stmt_33/bbx_xnph512_forx_xbody196_PhiReq/phi_stmt_677/phi_stmt_677_sources/$entry
      -- 
    ca_1314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_660_inst_ack_1, ack => convTranspose_CP_39_elements(168)); -- 
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	484 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	208 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_final_index_sum_regn_Sample/ack
      -- CP-element group 169: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_final_index_sum_regn_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_final_index_sum_regn_sample_complete
      -- 
    ack_1343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_689_index_offset_ack_0, ack => convTranspose_CP_39_elements(169)); -- 
    -- CP-element group 170:  transition  input  output  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	484 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	171 
    -- CP-element group 170:  members (11) 
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/addr_of_690_request/$entry
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_final_index_sum_regn_Update/ack
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_final_index_sum_regn_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/addr_of_690_request/req
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_base_plus_offset/sum_rename_ack
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_base_plus_offset/sum_rename_req
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_base_plus_offset/$exit
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_base_plus_offset/$entry
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_offset_calculated
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_root_address_calculated
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/addr_of_690_sample_start_
      -- 
    ack_1348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_689_index_offset_ack_1, ack => convTranspose_CP_39_elements(170)); -- 
    req_1357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(170), ack => addr_of_690_final_reg_req_0); -- 
    -- CP-element group 171:  transition  input  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	170 
    -- CP-element group 171: successors 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/addr_of_690_request/$exit
      -- CP-element group 171: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/addr_of_690_request/ack
      -- CP-element group 171: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/addr_of_690_sample_completed_
      -- 
    ack_1358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_690_final_reg_ack_0, ack => convTranspose_CP_39_elements(171)); -- 
    -- CP-element group 172:  fork  transition  input  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	484 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	205 
    -- CP-element group 172:  members (19) 
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/addr_of_690_complete/ack
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/addr_of_690_complete/$exit
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/addr_of_690_update_completed_
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_base_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_word_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_root_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_base_address_resized
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_base_addr_resize/$entry
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_base_addr_resize/$exit
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_base_addr_resize/base_resize_req
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_base_addr_resize/base_resize_ack
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_base_plus_offset/$entry
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_base_plus_offset/$exit
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_base_plus_offset/sum_rename_req
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_base_plus_offset/sum_rename_ack
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_word_addrgen/$entry
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_word_addrgen/$exit
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_word_addrgen/root_register_req
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_word_addrgen/root_register_ack
      -- 
    ack_1363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_690_final_reg_ack_1, ack => convTranspose_CP_39_elements(172)); -- 
    -- CP-element group 173:  transition  input  output  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	484 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	174 
    -- CP-element group 173:  members (6) 
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_693_Update/cr
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_693_Update/$entry
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_693_Sample/ra
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_693_Sample/$exit
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_693_update_start_
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_693_sample_completed_
      -- 
    ra_1372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_693_inst_ack_0, ack => convTranspose_CP_39_elements(173)); -- 
    cr_1376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(173), ack => RPIPE_ConvTranspose_input_pipe_693_inst_req_1); -- 
    -- CP-element group 174:  fork  transition  input  output  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	173 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	175 
    -- CP-element group 174: 	177 
    -- CP-element group 174:  members (9) 
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_706_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_697_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_706_Sample/rr
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_697_Sample/rr
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_697_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_706_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_693_Update/ca
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_693_Update/$exit
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_693_update_completed_
      -- 
    ca_1377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_693_inst_ack_1, ack => convTranspose_CP_39_elements(174)); -- 
    rr_1385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(174), ack => type_cast_697_inst_req_0); -- 
    rr_1399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(174), ack => RPIPE_ConvTranspose_input_pipe_706_inst_req_0); -- 
    -- CP-element group 175:  transition  input  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	174 
    -- CP-element group 175: successors 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_697_sample_completed_
      -- CP-element group 175: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_697_Sample/ra
      -- CP-element group 175: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_697_Sample/$exit
      -- 
    ra_1386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_697_inst_ack_0, ack => convTranspose_CP_39_elements(175)); -- 
    -- CP-element group 176:  transition  input  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	484 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	205 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_697_Update/ca
      -- CP-element group 176: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_697_Update/$exit
      -- CP-element group 176: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_697_update_completed_
      -- 
    ca_1391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_697_inst_ack_1, ack => convTranspose_CP_39_elements(176)); -- 
    -- CP-element group 177:  transition  input  output  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	174 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	178 
    -- CP-element group 177:  members (6) 
      -- CP-element group 177: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_706_sample_completed_
      -- CP-element group 177: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_706_Sample/ra
      -- CP-element group 177: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_706_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_706_Update/cr
      -- CP-element group 177: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_706_update_start_
      -- CP-element group 177: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_706_Update/$entry
      -- 
    ra_1400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_706_inst_ack_0, ack => convTranspose_CP_39_elements(177)); -- 
    cr_1404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(177), ack => RPIPE_ConvTranspose_input_pipe_706_inst_req_1); -- 
    -- CP-element group 178:  fork  transition  input  output  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	177 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178: 	181 
    -- CP-element group 178:  members (9) 
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_724_sample_start_
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_724_Sample/rr
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_724_Sample/$entry
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_706_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_706_Update/ca
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_710_sample_start_
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_710_Sample/rr
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_706_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_710_Sample/$entry
      -- 
    ca_1405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_706_inst_ack_1, ack => convTranspose_CP_39_elements(178)); -- 
    rr_1413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(178), ack => type_cast_710_inst_req_0); -- 
    rr_1427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(178), ack => RPIPE_ConvTranspose_input_pipe_724_inst_req_0); -- 
    -- CP-element group 179:  transition  input  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	178 
    -- CP-element group 179: successors 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_710_sample_completed_
      -- CP-element group 179: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_710_Sample/ra
      -- CP-element group 179: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_710_Sample/$exit
      -- 
    ra_1414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_710_inst_ack_0, ack => convTranspose_CP_39_elements(179)); -- 
    -- CP-element group 180:  transition  input  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	484 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	205 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_710_Update/ca
      -- CP-element group 180: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_710_Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_710_update_completed_
      -- 
    ca_1419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_710_inst_ack_1, ack => convTranspose_CP_39_elements(180)); -- 
    -- CP-element group 181:  transition  input  output  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	178 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	182 
    -- CP-element group 181:  members (6) 
      -- CP-element group 181: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_724_update_start_
      -- CP-element group 181: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_724_sample_completed_
      -- CP-element group 181: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_724_Sample/$exit
      -- CP-element group 181: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_724_Update/cr
      -- CP-element group 181: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_724_Update/$entry
      -- CP-element group 181: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_724_Sample/ra
      -- 
    ra_1428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_724_inst_ack_0, ack => convTranspose_CP_39_elements(181)); -- 
    cr_1432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(181), ack => RPIPE_ConvTranspose_input_pipe_724_inst_req_1); -- 
    -- CP-element group 182:  fork  transition  input  output  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	181 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	183 
    -- CP-element group 182: 	185 
    -- CP-element group 182:  members (9) 
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_728_Sample/rr
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_742_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_742_Sample/rr
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_742_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_724_update_completed_
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_728_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_728_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_724_Update/ca
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_724_Update/$exit
      -- 
    ca_1433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_724_inst_ack_1, ack => convTranspose_CP_39_elements(182)); -- 
    rr_1441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(182), ack => type_cast_728_inst_req_0); -- 
    rr_1455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(182), ack => RPIPE_ConvTranspose_input_pipe_742_inst_req_0); -- 
    -- CP-element group 183:  transition  input  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	182 
    -- CP-element group 183: successors 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_728_Sample/$exit
      -- CP-element group 183: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_728_Sample/ra
      -- CP-element group 183: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_728_sample_completed_
      -- 
    ra_1442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_728_inst_ack_0, ack => convTranspose_CP_39_elements(183)); -- 
    -- CP-element group 184:  transition  input  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	484 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	205 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_728_Update/ca
      -- CP-element group 184: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_728_update_completed_
      -- CP-element group 184: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_728_Update/$exit
      -- 
    ca_1447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_728_inst_ack_1, ack => convTranspose_CP_39_elements(184)); -- 
    -- CP-element group 185:  transition  input  output  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	182 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	186 
    -- CP-element group 185:  members (6) 
      -- CP-element group 185: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_742_Sample/$exit
      -- CP-element group 185: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_742_update_start_
      -- CP-element group 185: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_742_sample_completed_
      -- CP-element group 185: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_742_Sample/ra
      -- CP-element group 185: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_742_Update/$entry
      -- CP-element group 185: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_742_Update/cr
      -- 
    ra_1456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_742_inst_ack_0, ack => convTranspose_CP_39_elements(185)); -- 
    cr_1460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(185), ack => RPIPE_ConvTranspose_input_pipe_742_inst_req_1); -- 
    -- CP-element group 186:  fork  transition  input  output  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	185 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186: 	189 
    -- CP-element group 186:  members (9) 
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_742_update_completed_
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_742_Update/$exit
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_742_Update/ca
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_746_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_746_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_746_Sample/rr
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_760_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_760_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_760_Sample/rr
      -- 
    ca_1461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_742_inst_ack_1, ack => convTranspose_CP_39_elements(186)); -- 
    rr_1469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(186), ack => type_cast_746_inst_req_0); -- 
    rr_1483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(186), ack => RPIPE_ConvTranspose_input_pipe_760_inst_req_0); -- 
    -- CP-element group 187:  transition  input  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_746_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_746_Sample/$exit
      -- CP-element group 187: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_746_Sample/ra
      -- 
    ra_1470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_746_inst_ack_0, ack => convTranspose_CP_39_elements(187)); -- 
    -- CP-element group 188:  transition  input  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	484 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	205 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_746_update_completed_
      -- CP-element group 188: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_746_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_746_Update/ca
      -- 
    ca_1475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_746_inst_ack_1, ack => convTranspose_CP_39_elements(188)); -- 
    -- CP-element group 189:  transition  input  output  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	186 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	190 
    -- CP-element group 189:  members (6) 
      -- CP-element group 189: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_760_sample_completed_
      -- CP-element group 189: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_760_update_start_
      -- CP-element group 189: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_760_Sample/$exit
      -- CP-element group 189: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_760_Sample/ra
      -- CP-element group 189: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_760_Update/$entry
      -- CP-element group 189: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_760_Update/cr
      -- 
    ra_1484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_760_inst_ack_0, ack => convTranspose_CP_39_elements(189)); -- 
    cr_1488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(189), ack => RPIPE_ConvTranspose_input_pipe_760_inst_req_1); -- 
    -- CP-element group 190:  fork  transition  input  output  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	189 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	191 
    -- CP-element group 190: 	193 
    -- CP-element group 190:  members (9) 
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_760_update_completed_
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_760_Update/$exit
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_760_Update/ca
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_764_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_764_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_764_Sample/rr
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_778_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_778_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_778_Sample/rr
      -- 
    ca_1489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_760_inst_ack_1, ack => convTranspose_CP_39_elements(190)); -- 
    rr_1497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(190), ack => type_cast_764_inst_req_0); -- 
    rr_1511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(190), ack => RPIPE_ConvTranspose_input_pipe_778_inst_req_0); -- 
    -- CP-element group 191:  transition  input  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	190 
    -- CP-element group 191: successors 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_764_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_764_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_764_Sample/ra
      -- 
    ra_1498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_764_inst_ack_0, ack => convTranspose_CP_39_elements(191)); -- 
    -- CP-element group 192:  transition  input  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	484 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	205 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_764_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_764_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_764_Update/ca
      -- 
    ca_1503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_764_inst_ack_1, ack => convTranspose_CP_39_elements(192)); -- 
    -- CP-element group 193:  transition  input  output  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	190 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	194 
    -- CP-element group 193:  members (6) 
      -- CP-element group 193: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_778_sample_completed_
      -- CP-element group 193: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_778_update_start_
      -- CP-element group 193: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_778_Sample/$exit
      -- CP-element group 193: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_778_Sample/ra
      -- CP-element group 193: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_778_Update/$entry
      -- CP-element group 193: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_778_Update/cr
      -- 
    ra_1512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_778_inst_ack_0, ack => convTranspose_CP_39_elements(193)); -- 
    cr_1516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(193), ack => RPIPE_ConvTranspose_input_pipe_778_inst_req_1); -- 
    -- CP-element group 194:  fork  transition  input  output  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	193 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194: 	197 
    -- CP-element group 194:  members (9) 
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_778_update_completed_
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_778_Update/$exit
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_778_Update/ca
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_782_sample_start_
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_782_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_782_Sample/rr
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_796_sample_start_
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_796_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_796_Sample/rr
      -- 
    ca_1517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_778_inst_ack_1, ack => convTranspose_CP_39_elements(194)); -- 
    rr_1525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(194), ack => type_cast_782_inst_req_0); -- 
    rr_1539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(194), ack => RPIPE_ConvTranspose_input_pipe_796_inst_req_0); -- 
    -- CP-element group 195:  transition  input  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_782_sample_completed_
      -- CP-element group 195: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_782_Sample/$exit
      -- CP-element group 195: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_782_Sample/ra
      -- 
    ra_1526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_782_inst_ack_0, ack => convTranspose_CP_39_elements(195)); -- 
    -- CP-element group 196:  transition  input  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	484 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	205 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_782_update_completed_
      -- CP-element group 196: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_782_Update/$exit
      -- CP-element group 196: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_782_Update/ca
      -- 
    ca_1531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_782_inst_ack_1, ack => convTranspose_CP_39_elements(196)); -- 
    -- CP-element group 197:  transition  input  output  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	194 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	198 
    -- CP-element group 197:  members (6) 
      -- CP-element group 197: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_796_sample_completed_
      -- CP-element group 197: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_796_update_start_
      -- CP-element group 197: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_796_Sample/$exit
      -- CP-element group 197: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_796_Sample/ra
      -- CP-element group 197: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_796_Update/$entry
      -- CP-element group 197: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_796_Update/cr
      -- 
    ra_1540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_796_inst_ack_0, ack => convTranspose_CP_39_elements(197)); -- 
    cr_1544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(197), ack => RPIPE_ConvTranspose_input_pipe_796_inst_req_1); -- 
    -- CP-element group 198:  fork  transition  input  output  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	197 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	199 
    -- CP-element group 198: 	201 
    -- CP-element group 198:  members (9) 
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_796_update_completed_
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_796_Update/$exit
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_796_Update/ca
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_800_sample_start_
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_800_Sample/$entry
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_800_Sample/rr
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_814_sample_start_
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_814_Sample/$entry
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_814_Sample/rr
      -- 
    ca_1545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_796_inst_ack_1, ack => convTranspose_CP_39_elements(198)); -- 
    rr_1553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(198), ack => type_cast_800_inst_req_0); -- 
    rr_1567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(198), ack => RPIPE_ConvTranspose_input_pipe_814_inst_req_0); -- 
    -- CP-element group 199:  transition  input  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	198 
    -- CP-element group 199: successors 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_800_sample_completed_
      -- CP-element group 199: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_800_Sample/$exit
      -- CP-element group 199: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_800_Sample/ra
      -- 
    ra_1554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_800_inst_ack_0, ack => convTranspose_CP_39_elements(199)); -- 
    -- CP-element group 200:  transition  input  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	484 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	205 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_800_update_completed_
      -- CP-element group 200: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_800_Update/$exit
      -- CP-element group 200: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_800_Update/ca
      -- 
    ca_1559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_800_inst_ack_1, ack => convTranspose_CP_39_elements(200)); -- 
    -- CP-element group 201:  transition  input  output  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	198 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201:  members (6) 
      -- CP-element group 201: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_814_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_814_update_start_
      -- CP-element group 201: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_814_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_814_Sample/ra
      -- CP-element group 201: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_814_Update/$entry
      -- CP-element group 201: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_814_Update/cr
      -- 
    ra_1568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_814_inst_ack_0, ack => convTranspose_CP_39_elements(201)); -- 
    cr_1572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(201), ack => RPIPE_ConvTranspose_input_pipe_814_inst_req_1); -- 
    -- CP-element group 202:  transition  input  output  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	201 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202:  members (6) 
      -- CP-element group 202: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_814_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_814_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_814_Update/ca
      -- CP-element group 202: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_818_sample_start_
      -- CP-element group 202: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_818_Sample/$entry
      -- CP-element group 202: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_818_Sample/rr
      -- 
    ca_1573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_814_inst_ack_1, ack => convTranspose_CP_39_elements(202)); -- 
    rr_1581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(202), ack => type_cast_818_inst_req_0); -- 
    -- CP-element group 203:  transition  input  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	202 
    -- CP-element group 203: successors 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_818_sample_completed_
      -- CP-element group 203: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_818_Sample/$exit
      -- CP-element group 203: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_818_Sample/ra
      -- 
    ra_1582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_818_inst_ack_0, ack => convTranspose_CP_39_elements(203)); -- 
    -- CP-element group 204:  transition  input  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	484 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	205 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_818_update_completed_
      -- CP-element group 204: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_818_Update/$exit
      -- CP-element group 204: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_818_Update/ca
      -- 
    ca_1587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_818_inst_ack_1, ack => convTranspose_CP_39_elements(204)); -- 
    -- CP-element group 205:  join  transition  output  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	180 
    -- CP-element group 205: 	184 
    -- CP-element group 205: 	188 
    -- CP-element group 205: 	192 
    -- CP-element group 205: 	196 
    -- CP-element group 205: 	200 
    -- CP-element group 205: 	204 
    -- CP-element group 205: 	176 
    -- CP-element group 205: 	172 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	206 
    -- CP-element group 205:  members (9) 
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_sample_start_
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_Sample/$entry
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_Sample/ptr_deref_826_Split/$entry
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_Sample/ptr_deref_826_Split/$exit
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_Sample/ptr_deref_826_Split/split_req
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_Sample/ptr_deref_826_Split/split_ack
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_Sample/word_access_start/$entry
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_Sample/word_access_start/word_0/$entry
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_Sample/word_access_start/word_0/rr
      -- 
    rr_1625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(205), ack => ptr_deref_826_store_0_req_0); -- 
    convTranspose_cp_element_group_205: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_205"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(180) & convTranspose_CP_39_elements(184) & convTranspose_CP_39_elements(188) & convTranspose_CP_39_elements(192) & convTranspose_CP_39_elements(196) & convTranspose_CP_39_elements(200) & convTranspose_CP_39_elements(204) & convTranspose_CP_39_elements(176) & convTranspose_CP_39_elements(172);
      gj_convTranspose_cp_element_group_205 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(205), clk => clk, reset => reset); --
    end block;
    -- CP-element group 206:  transition  input  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	205 
    -- CP-element group 206: successors 
    -- CP-element group 206:  members (5) 
      -- CP-element group 206: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_sample_completed_
      -- CP-element group 206: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_Sample/$exit
      -- CP-element group 206: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_Sample/word_access_start/$exit
      -- CP-element group 206: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_Sample/word_access_start/word_0/$exit
      -- CP-element group 206: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_Sample/word_access_start/word_0/ra
      -- 
    ra_1626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_826_store_0_ack_0, ack => convTranspose_CP_39_elements(206)); -- 
    -- CP-element group 207:  transition  input  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	484 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	208 
    -- CP-element group 207:  members (5) 
      -- CP-element group 207: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_update_completed_
      -- CP-element group 207: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_Update/$exit
      -- CP-element group 207: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_Update/word_access_complete/$exit
      -- CP-element group 207: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_Update/word_access_complete/word_0/$exit
      -- CP-element group 207: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_Update/word_access_complete/word_0/ca
      -- 
    ca_1637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_826_store_0_ack_1, ack => convTranspose_CP_39_elements(207)); -- 
    -- CP-element group 208:  branch  join  transition  place  output  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	207 
    -- CP-element group 208: 	169 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	209 
    -- CP-element group 208: 	210 
    -- CP-element group 208:  members (10) 
      -- CP-element group 208: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839__exit__
      -- CP-element group 208: 	 branch_block_stmt_33/if_stmt_840__entry__
      -- CP-element group 208: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/$exit
      -- CP-element group 208: 	 branch_block_stmt_33/if_stmt_840_dead_link/$entry
      -- CP-element group 208: 	 branch_block_stmt_33/if_stmt_840_eval_test/$entry
      -- CP-element group 208: 	 branch_block_stmt_33/if_stmt_840_eval_test/$exit
      -- CP-element group 208: 	 branch_block_stmt_33/if_stmt_840_eval_test/branch_req
      -- CP-element group 208: 	 branch_block_stmt_33/R_exitcond2_841_place
      -- CP-element group 208: 	 branch_block_stmt_33/if_stmt_840_if_link/$entry
      -- CP-element group 208: 	 branch_block_stmt_33/if_stmt_840_else_link/$entry
      -- 
    branch_req_1645_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1645_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(208), ack => if_stmt_840_branch_req_0); -- 
    convTranspose_cp_element_group_208: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_208"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(207) & convTranspose_CP_39_elements(169);
      gj_convTranspose_cp_element_group_208 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(208), clk => clk, reset => reset); --
    end block;
    -- CP-element group 209:  merge  transition  place  input  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	208 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	485 
    -- CP-element group 209:  members (13) 
      -- CP-element group 209: 	 branch_block_stmt_33/merge_stmt_846__exit__
      -- CP-element group 209: 	 branch_block_stmt_33/forx_xend250x_xloopexit_forx_xend250
      -- CP-element group 209: 	 branch_block_stmt_33/if_stmt_840_if_link/$exit
      -- CP-element group 209: 	 branch_block_stmt_33/if_stmt_840_if_link/if_choice_transition
      -- CP-element group 209: 	 branch_block_stmt_33/forx_xbody196_forx_xend250x_xloopexit
      -- CP-element group 209: 	 branch_block_stmt_33/forx_xbody196_forx_xend250x_xloopexit_PhiReq/$entry
      -- CP-element group 209: 	 branch_block_stmt_33/forx_xbody196_forx_xend250x_xloopexit_PhiReq/$exit
      -- CP-element group 209: 	 branch_block_stmt_33/merge_stmt_846_PhiReqMerge
      -- CP-element group 209: 	 branch_block_stmt_33/merge_stmt_846_PhiAck/$entry
      -- CP-element group 209: 	 branch_block_stmt_33/merge_stmt_846_PhiAck/$exit
      -- CP-element group 209: 	 branch_block_stmt_33/merge_stmt_846_PhiAck/dummy
      -- CP-element group 209: 	 branch_block_stmt_33/forx_xend250x_xloopexit_forx_xend250_PhiReq/$entry
      -- CP-element group 209: 	 branch_block_stmt_33/forx_xend250x_xloopexit_forx_xend250_PhiReq/$exit
      -- 
    if_choice_transition_1650_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_840_branch_ack_1, ack => convTranspose_CP_39_elements(209)); -- 
    -- CP-element group 210:  fork  transition  place  input  output  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	208 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	480 
    -- CP-element group 210: 	481 
    -- CP-element group 210:  members (12) 
      -- CP-element group 210: 	 branch_block_stmt_33/if_stmt_840_else_link/$exit
      -- CP-element group 210: 	 branch_block_stmt_33/if_stmt_840_else_link/else_choice_transition
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody196_forx_xbody196
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody196_forx_xbody196_PhiReq/$entry
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_677/$entry
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_677/phi_stmt_677_sources/$entry
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_677/phi_stmt_677_sources/type_cast_683/$entry
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_677/phi_stmt_677_sources/type_cast_683/SplitProtocol/$entry
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_677/phi_stmt_677_sources/type_cast_683/SplitProtocol/Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_677/phi_stmt_677_sources/type_cast_683/SplitProtocol/Sample/rr
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_677/phi_stmt_677_sources/type_cast_683/SplitProtocol/Update/$entry
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_677/phi_stmt_677_sources/type_cast_683/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_840_branch_ack_0, ack => convTranspose_CP_39_elements(210)); -- 
    rr_3579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(210), ack => type_cast_683_inst_req_0); -- 
    cr_3584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(210), ack => type_cast_683_inst_req_1); -- 
    -- CP-element group 211:  transition  input  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	485 
    -- CP-element group 211: successors 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_851_sample_completed_
      -- CP-element group 211: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_851_Sample/$exit
      -- CP-element group 211: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_851_Sample/ra
      -- 
    ra_1668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_851_inst_ack_0, ack => convTranspose_CP_39_elements(211)); -- 
    -- CP-element group 212:  transition  input  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	485 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	217 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_851_update_completed_
      -- CP-element group 212: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_851_Update/$exit
      -- CP-element group 212: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_851_Update/ca
      -- 
    ca_1673_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_851_inst_ack_1, ack => convTranspose_CP_39_elements(212)); -- 
    -- CP-element group 213:  transition  input  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	485 
    -- CP-element group 213: successors 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_855_sample_completed_
      -- CP-element group 213: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_855_Sample/$exit
      -- CP-element group 213: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_855_Sample/ra
      -- 
    ra_1682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_855_inst_ack_0, ack => convTranspose_CP_39_elements(213)); -- 
    -- CP-element group 214:  transition  input  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	485 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	217 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_855_update_completed_
      -- CP-element group 214: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_855_Update/$exit
      -- CP-element group 214: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_855_Update/ca
      -- 
    ca_1687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_855_inst_ack_1, ack => convTranspose_CP_39_elements(214)); -- 
    -- CP-element group 215:  transition  input  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	485 
    -- CP-element group 215: successors 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_859_sample_completed_
      -- CP-element group 215: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_859_Sample/$exit
      -- CP-element group 215: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_859_Sample/ra
      -- 
    ra_1696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_859_inst_ack_0, ack => convTranspose_CP_39_elements(215)); -- 
    -- CP-element group 216:  transition  input  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	485 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	217 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_859_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_859_Update/$exit
      -- CP-element group 216: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_859_Update/ca
      -- 
    ca_1701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_859_inst_ack_1, ack => convTranspose_CP_39_elements(216)); -- 
    -- CP-element group 217:  branch  join  transition  place  output  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	212 
    -- CP-element group 217: 	214 
    -- CP-element group 217: 	216 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	218 
    -- CP-element group 217: 	219 
    -- CP-element group 217:  members (10) 
      -- CP-element group 217: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876__exit__
      -- CP-element group 217: 	 branch_block_stmt_33/if_stmt_877__entry__
      -- CP-element group 217: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/$exit
      -- CP-element group 217: 	 branch_block_stmt_33/if_stmt_877_dead_link/$entry
      -- CP-element group 217: 	 branch_block_stmt_33/if_stmt_877_eval_test/$entry
      -- CP-element group 217: 	 branch_block_stmt_33/if_stmt_877_eval_test/$exit
      -- CP-element group 217: 	 branch_block_stmt_33/if_stmt_877_eval_test/branch_req
      -- CP-element group 217: 	 branch_block_stmt_33/R_cmp264506_878_place
      -- CP-element group 217: 	 branch_block_stmt_33/if_stmt_877_if_link/$entry
      -- CP-element group 217: 	 branch_block_stmt_33/if_stmt_877_else_link/$entry
      -- 
    branch_req_1709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(217), ack => if_stmt_877_branch_req_0); -- 
    convTranspose_cp_element_group_217: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_217"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(212) & convTranspose_CP_39_elements(214) & convTranspose_CP_39_elements(216);
      gj_convTranspose_cp_element_group_217 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(217), clk => clk, reset => reset); --
    end block;
    -- CP-element group 218:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	217 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	220 
    -- CP-element group 218: 	221 
    -- CP-element group 218:  members (18) 
      -- CP-element group 218: 	 branch_block_stmt_33/merge_stmt_883__exit__
      -- CP-element group 218: 	 branch_block_stmt_33/assign_stmt_889_to_assign_stmt_918__entry__
      -- CP-element group 218: 	 branch_block_stmt_33/if_stmt_877_if_link/$exit
      -- CP-element group 218: 	 branch_block_stmt_33/if_stmt_877_if_link/if_choice_transition
      -- CP-element group 218: 	 branch_block_stmt_33/forx_xend250_bbx_xnph508
      -- CP-element group 218: 	 branch_block_stmt_33/assign_stmt_889_to_assign_stmt_918/$entry
      -- CP-element group 218: 	 branch_block_stmt_33/assign_stmt_889_to_assign_stmt_918/type_cast_904_sample_start_
      -- CP-element group 218: 	 branch_block_stmt_33/assign_stmt_889_to_assign_stmt_918/type_cast_904_update_start_
      -- CP-element group 218: 	 branch_block_stmt_33/assign_stmt_889_to_assign_stmt_918/type_cast_904_Sample/$entry
      -- CP-element group 218: 	 branch_block_stmt_33/assign_stmt_889_to_assign_stmt_918/type_cast_904_Sample/rr
      -- CP-element group 218: 	 branch_block_stmt_33/assign_stmt_889_to_assign_stmt_918/type_cast_904_Update/$entry
      -- CP-element group 218: 	 branch_block_stmt_33/assign_stmt_889_to_assign_stmt_918/type_cast_904_Update/cr
      -- CP-element group 218: 	 branch_block_stmt_33/forx_xend250_bbx_xnph508_PhiReq/$entry
      -- CP-element group 218: 	 branch_block_stmt_33/forx_xend250_bbx_xnph508_PhiReq/$exit
      -- CP-element group 218: 	 branch_block_stmt_33/merge_stmt_883_PhiReqMerge
      -- CP-element group 218: 	 branch_block_stmt_33/merge_stmt_883_PhiAck/$entry
      -- CP-element group 218: 	 branch_block_stmt_33/merge_stmt_883_PhiAck/$exit
      -- CP-element group 218: 	 branch_block_stmt_33/merge_stmt_883_PhiAck/dummy
      -- 
    if_choice_transition_1714_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_877_branch_ack_1, ack => convTranspose_CP_39_elements(218)); -- 
    rr_1731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(218), ack => type_cast_904_inst_req_0); -- 
    cr_1736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(218), ack => type_cast_904_inst_req_1); -- 
    -- CP-element group 219:  transition  place  input  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	217 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	492 
    -- CP-element group 219:  members (5) 
      -- CP-element group 219: 	 branch_block_stmt_33/if_stmt_877_else_link/$exit
      -- CP-element group 219: 	 branch_block_stmt_33/if_stmt_877_else_link/else_choice_transition
      -- CP-element group 219: 	 branch_block_stmt_33/forx_xend250_forx_xend273
      -- CP-element group 219: 	 branch_block_stmt_33/forx_xend250_forx_xend273_PhiReq/$entry
      -- CP-element group 219: 	 branch_block_stmt_33/forx_xend250_forx_xend273_PhiReq/$exit
      -- 
    else_choice_transition_1718_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_877_branch_ack_0, ack => convTranspose_CP_39_elements(219)); -- 
    -- CP-element group 220:  transition  input  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	218 
    -- CP-element group 220: successors 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_33/assign_stmt_889_to_assign_stmt_918/type_cast_904_sample_completed_
      -- CP-element group 220: 	 branch_block_stmt_33/assign_stmt_889_to_assign_stmt_918/type_cast_904_Sample/$exit
      -- CP-element group 220: 	 branch_block_stmt_33/assign_stmt_889_to_assign_stmt_918/type_cast_904_Sample/ra
      -- 
    ra_1732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_904_inst_ack_0, ack => convTranspose_CP_39_elements(220)); -- 
    -- CP-element group 221:  transition  place  input  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	218 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	486 
    -- CP-element group 221:  members (9) 
      -- CP-element group 221: 	 branch_block_stmt_33/assign_stmt_889_to_assign_stmt_918__exit__
      -- CP-element group 221: 	 branch_block_stmt_33/bbx_xnph508_forx_xbody266
      -- CP-element group 221: 	 branch_block_stmt_33/assign_stmt_889_to_assign_stmt_918/$exit
      -- CP-element group 221: 	 branch_block_stmt_33/assign_stmt_889_to_assign_stmt_918/type_cast_904_update_completed_
      -- CP-element group 221: 	 branch_block_stmt_33/assign_stmt_889_to_assign_stmt_918/type_cast_904_Update/$exit
      -- CP-element group 221: 	 branch_block_stmt_33/assign_stmt_889_to_assign_stmt_918/type_cast_904_Update/ca
      -- CP-element group 221: 	 branch_block_stmt_33/bbx_xnph508_forx_xbody266_PhiReq/$entry
      -- CP-element group 221: 	 branch_block_stmt_33/bbx_xnph508_forx_xbody266_PhiReq/phi_stmt_921/$entry
      -- CP-element group 221: 	 branch_block_stmt_33/bbx_xnph508_forx_xbody266_PhiReq/phi_stmt_921/phi_stmt_921_sources/$entry
      -- 
    ca_1737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_904_inst_ack_1, ack => convTranspose_CP_39_elements(221)); -- 
    -- CP-element group 222:  transition  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	491 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	228 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_final_index_sum_regn_sample_complete
      -- CP-element group 222: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_final_index_sum_regn_Sample/$exit
      -- CP-element group 222: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_final_index_sum_regn_Sample/ack
      -- 
    ack_1766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_933_index_offset_ack_0, ack => convTranspose_CP_39_elements(222)); -- 
    -- CP-element group 223:  transition  input  output  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	491 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223:  members (11) 
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/addr_of_934_sample_start_
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_root_address_calculated
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_offset_calculated
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_final_index_sum_regn_Update/$exit
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_final_index_sum_regn_Update/ack
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_base_plus_offset/$entry
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_base_plus_offset/$exit
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_base_plus_offset/sum_rename_req
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_base_plus_offset/sum_rename_ack
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/addr_of_934_request/$entry
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/addr_of_934_request/req
      -- 
    ack_1771_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_933_index_offset_ack_1, ack => convTranspose_CP_39_elements(223)); -- 
    req_1780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(223), ack => addr_of_934_final_reg_req_0); -- 
    -- CP-element group 224:  transition  input  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/addr_of_934_sample_completed_
      -- CP-element group 224: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/addr_of_934_request/$exit
      -- CP-element group 224: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/addr_of_934_request/ack
      -- 
    ack_1781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_934_final_reg_ack_0, ack => convTranspose_CP_39_elements(224)); -- 
    -- CP-element group 225:  join  fork  transition  input  output  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	491 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	226 
    -- CP-element group 225:  members (28) 
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/addr_of_934_update_completed_
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/addr_of_934_complete/$exit
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/addr_of_934_complete/ack
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_sample_start_
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_base_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_word_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_root_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_base_address_resized
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_base_addr_resize/$entry
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_base_addr_resize/$exit
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_base_addr_resize/base_resize_req
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_base_addr_resize/base_resize_ack
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_base_plus_offset/$entry
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_base_plus_offset/$exit
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_base_plus_offset/sum_rename_req
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_base_plus_offset/sum_rename_ack
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_word_addrgen/$entry
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_word_addrgen/$exit
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_word_addrgen/root_register_req
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_word_addrgen/root_register_ack
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_Sample/$entry
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_Sample/ptr_deref_937_Split/$entry
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_Sample/ptr_deref_937_Split/$exit
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_Sample/ptr_deref_937_Split/split_req
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_Sample/ptr_deref_937_Split/split_ack
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_Sample/word_access_start/$entry
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_Sample/word_access_start/word_0/$entry
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_Sample/word_access_start/word_0/rr
      -- 
    ack_1786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_934_final_reg_ack_1, ack => convTranspose_CP_39_elements(225)); -- 
    rr_1824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(225), ack => ptr_deref_937_store_0_req_0); -- 
    -- CP-element group 226:  transition  input  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	225 
    -- CP-element group 226: successors 
    -- CP-element group 226:  members (5) 
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_sample_completed_
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_Sample/$exit
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_Sample/word_access_start/$exit
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_Sample/word_access_start/word_0/$exit
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_Sample/word_access_start/word_0/ra
      -- 
    ra_1825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_937_store_0_ack_0, ack => convTranspose_CP_39_elements(226)); -- 
    -- CP-element group 227:  transition  input  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	491 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	228 
    -- CP-element group 227:  members (5) 
      -- CP-element group 227: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_update_completed_
      -- CP-element group 227: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_Update/$exit
      -- CP-element group 227: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_Update/word_access_complete/$exit
      -- CP-element group 227: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_Update/word_access_complete/word_0/$exit
      -- CP-element group 227: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_Update/word_access_complete/word_0/ca
      -- 
    ca_1836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_937_store_0_ack_1, ack => convTranspose_CP_39_elements(227)); -- 
    -- CP-element group 228:  branch  join  transition  place  output  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	222 
    -- CP-element group 228: 	227 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	229 
    -- CP-element group 228: 	230 
    -- CP-element group 228:  members (10) 
      -- CP-element group 228: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951__exit__
      -- CP-element group 228: 	 branch_block_stmt_33/if_stmt_952__entry__
      -- CP-element group 228: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/$exit
      -- CP-element group 228: 	 branch_block_stmt_33/if_stmt_952_dead_link/$entry
      -- CP-element group 228: 	 branch_block_stmt_33/if_stmt_952_eval_test/$entry
      -- CP-element group 228: 	 branch_block_stmt_33/if_stmt_952_eval_test/$exit
      -- CP-element group 228: 	 branch_block_stmt_33/if_stmt_952_eval_test/branch_req
      -- CP-element group 228: 	 branch_block_stmt_33/R_exitcond_953_place
      -- CP-element group 228: 	 branch_block_stmt_33/if_stmt_952_if_link/$entry
      -- CP-element group 228: 	 branch_block_stmt_33/if_stmt_952_else_link/$entry
      -- 
    branch_req_1844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(228), ack => if_stmt_952_branch_req_0); -- 
    convTranspose_cp_element_group_228: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_228"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(222) & convTranspose_CP_39_elements(227);
      gj_convTranspose_cp_element_group_228 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(228), clk => clk, reset => reset); --
    end block;
    -- CP-element group 229:  merge  transition  place  input  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	228 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	492 
    -- CP-element group 229:  members (13) 
      -- CP-element group 229: 	 branch_block_stmt_33/merge_stmt_958__exit__
      -- CP-element group 229: 	 branch_block_stmt_33/forx_xend273x_xloopexit_forx_xend273
      -- CP-element group 229: 	 branch_block_stmt_33/if_stmt_952_if_link/$exit
      -- CP-element group 229: 	 branch_block_stmt_33/if_stmt_952_if_link/if_choice_transition
      -- CP-element group 229: 	 branch_block_stmt_33/forx_xbody266_forx_xend273x_xloopexit
      -- CP-element group 229: 	 branch_block_stmt_33/forx_xbody266_forx_xend273x_xloopexit_PhiReq/$entry
      -- CP-element group 229: 	 branch_block_stmt_33/forx_xbody266_forx_xend273x_xloopexit_PhiReq/$exit
      -- CP-element group 229: 	 branch_block_stmt_33/merge_stmt_958_PhiReqMerge
      -- CP-element group 229: 	 branch_block_stmt_33/merge_stmt_958_PhiAck/$entry
      -- CP-element group 229: 	 branch_block_stmt_33/merge_stmt_958_PhiAck/$exit
      -- CP-element group 229: 	 branch_block_stmt_33/merge_stmt_958_PhiAck/dummy
      -- CP-element group 229: 	 branch_block_stmt_33/forx_xend273x_xloopexit_forx_xend273_PhiReq/$entry
      -- CP-element group 229: 	 branch_block_stmt_33/forx_xend273x_xloopexit_forx_xend273_PhiReq/$exit
      -- 
    if_choice_transition_1849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_952_branch_ack_1, ack => convTranspose_CP_39_elements(229)); -- 
    -- CP-element group 230:  fork  transition  place  input  output  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	228 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	487 
    -- CP-element group 230: 	488 
    -- CP-element group 230:  members (12) 
      -- CP-element group 230: 	 branch_block_stmt_33/if_stmt_952_else_link/$exit
      -- CP-element group 230: 	 branch_block_stmt_33/if_stmt_952_else_link/else_choice_transition
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody266_forx_xbody266
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody266_forx_xbody266_PhiReq/$entry
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_921/$entry
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_921/phi_stmt_921_sources/$entry
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_921/phi_stmt_921_sources/type_cast_924/$entry
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_921/phi_stmt_921_sources/type_cast_924/SplitProtocol/$entry
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_921/phi_stmt_921_sources/type_cast_924/SplitProtocol/Sample/$entry
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_921/phi_stmt_921_sources/type_cast_924/SplitProtocol/Sample/rr
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_921/phi_stmt_921_sources/type_cast_924/SplitProtocol/Update/$entry
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_921/phi_stmt_921_sources/type_cast_924/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_952_branch_ack_0, ack => convTranspose_CP_39_elements(230)); -- 
    rr_3656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(230), ack => type_cast_924_inst_req_0); -- 
    cr_3661_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3661_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(230), ack => type_cast_924_inst_req_1); -- 
    -- CP-element group 231:  transition  input  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	492 
    -- CP-element group 231: successors 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_969/call_stmt_963_sample_completed_
      -- CP-element group 231: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_969/call_stmt_963_Sample/$exit
      -- CP-element group 231: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_969/call_stmt_963_Sample/cra
      -- 
    cra_1867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_963_call_ack_0, ack => convTranspose_CP_39_elements(231)); -- 
    -- CP-element group 232:  transition  input  output  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	492 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	233 
    -- CP-element group 232:  members (6) 
      -- CP-element group 232: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_969/call_stmt_963_update_completed_
      -- CP-element group 232: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_969/call_stmt_963_Update/$exit
      -- CP-element group 232: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_969/call_stmt_963_Update/cca
      -- CP-element group 232: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_969/type_cast_968_sample_start_
      -- CP-element group 232: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_969/type_cast_968_Sample/$entry
      -- CP-element group 232: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_969/type_cast_968_Sample/rr
      -- 
    cca_1872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_963_call_ack_1, ack => convTranspose_CP_39_elements(232)); -- 
    rr_1880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(232), ack => type_cast_968_inst_req_0); -- 
    -- CP-element group 233:  transition  input  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	232 
    -- CP-element group 233: successors 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_969/type_cast_968_sample_completed_
      -- CP-element group 233: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_969/type_cast_968_Sample/$exit
      -- CP-element group 233: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_969/type_cast_968_Sample/ra
      -- 
    ra_1881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_968_inst_ack_0, ack => convTranspose_CP_39_elements(233)); -- 
    -- CP-element group 234:  fork  transition  place  input  output  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	492 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	331 
    -- CP-element group 234: 	349 
    -- CP-element group 234: 	350 
    -- CP-element group 234: 	354 
    -- CP-element group 234: 	355 
    -- CP-element group 234: 	365 
    -- CP-element group 234: 	367 
    -- CP-element group 234: 	369 
    -- CP-element group 234: 	371 
    -- CP-element group 234: 	235 
    -- CP-element group 234: 	263 
    -- CP-element group 234: 	281 
    -- CP-element group 234: 	282 
    -- CP-element group 234: 	286 
    -- CP-element group 234: 	287 
    -- CP-element group 234: 	297 
    -- CP-element group 234: 	315 
    -- CP-element group 234: 	316 
    -- CP-element group 234: 	320 
    -- CP-element group 234: 	321 
    -- CP-element group 234:  members (67) 
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1071_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1106_update_start_
      -- CP-element group 234: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_969__exit__
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194__entry__
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1050_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1050_update_start_
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1071_Sample/req
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1050_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1050_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1050_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1071_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1050_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1057_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1057_update_start_
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1057_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1057_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1057_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1106_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1015_Sample/req
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1015_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1015_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1057_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_969/$exit
      -- CP-element group 234: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_969/type_cast_968_update_completed_
      -- CP-element group 234: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_969/type_cast_968_Update/$exit
      -- CP-element group 234: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_969/type_cast_968_Update/ca
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/$entry
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_971_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_971_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_971_Sample/req
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1106_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1106_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1106_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1106_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1113_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1113_update_start_
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1113_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1113_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1113_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1113_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1127_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1127_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1127_Sample/req
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1162_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1162_update_start_
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1162_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1162_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1162_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1162_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1169_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1169_update_start_
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1169_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1169_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1169_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1169_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block0_done_1184_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block0_done_1184_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block0_done_1184_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block1_done_1187_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block1_done_1187_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block1_done_1187_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block2_done_1190_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block2_done_1190_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block2_done_1190_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block3_done_1193_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block3_done_1193_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block3_done_1193_Sample/rr
      -- 
    ca_1886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_968_inst_ack_1, ack => convTranspose_CP_39_elements(234)); -- 
    req_2317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => WPIPE_Block2_start_1071_inst_req_0); -- 
    cr_2224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => type_cast_1050_inst_req_1); -- 
    rr_2219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => type_cast_1050_inst_req_0); -- 
    rr_2247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => type_cast_1057_inst_req_0); -- 
    req_2093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => WPIPE_Block1_start_1015_inst_req_0); -- 
    cr_2252_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2252_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => type_cast_1057_inst_req_1); -- 
    req_1897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => WPIPE_Block0_start_971_inst_req_0); -- 
    rr_2443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => type_cast_1106_inst_req_0); -- 
    cr_2448_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2448_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => type_cast_1106_inst_req_1); -- 
    rr_2471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => type_cast_1113_inst_req_0); -- 
    cr_2476_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2476_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => type_cast_1113_inst_req_1); -- 
    req_2541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => WPIPE_Block3_start_1127_inst_req_0); -- 
    rr_2667_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2667_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => type_cast_1162_inst_req_0); -- 
    cr_2672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => type_cast_1162_inst_req_1); -- 
    rr_2695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => type_cast_1169_inst_req_0); -- 
    cr_2700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => type_cast_1169_inst_req_1); -- 
    rr_2765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => RPIPE_Block0_done_1184_inst_req_0); -- 
    rr_2779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => RPIPE_Block1_done_1187_inst_req_0); -- 
    rr_2793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => RPIPE_Block2_done_1190_inst_req_0); -- 
    rr_2807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => RPIPE_Block3_done_1193_inst_req_0); -- 
    -- CP-element group 235:  transition  input  output  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	234 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235:  members (6) 
      -- CP-element group 235: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_971_sample_completed_
      -- CP-element group 235: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_971_update_start_
      -- CP-element group 235: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_971_Sample/$exit
      -- CP-element group 235: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_971_Sample/ack
      -- CP-element group 235: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_971_Update/$entry
      -- CP-element group 235: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_971_Update/req
      -- 
    ack_1898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_971_inst_ack_0, ack => convTranspose_CP_39_elements(235)); -- 
    req_1902_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1902_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(235), ack => WPIPE_Block0_start_971_inst_req_1); -- 
    -- CP-element group 236:  transition  input  output  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	237 
    -- CP-element group 236:  members (6) 
      -- CP-element group 236: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_971_update_completed_
      -- CP-element group 236: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_971_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_971_Update/ack
      -- CP-element group 236: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_974_sample_start_
      -- CP-element group 236: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_974_Sample/$entry
      -- CP-element group 236: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_974_Sample/req
      -- 
    ack_1903_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_971_inst_ack_1, ack => convTranspose_CP_39_elements(236)); -- 
    req_1911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(236), ack => WPIPE_Block0_start_974_inst_req_0); -- 
    -- CP-element group 237:  transition  input  output  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	236 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	238 
    -- CP-element group 237:  members (6) 
      -- CP-element group 237: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_974_sample_completed_
      -- CP-element group 237: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_974_update_start_
      -- CP-element group 237: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_974_Sample/$exit
      -- CP-element group 237: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_974_Sample/ack
      -- CP-element group 237: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_974_Update/$entry
      -- CP-element group 237: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_974_Update/req
      -- 
    ack_1912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_974_inst_ack_0, ack => convTranspose_CP_39_elements(237)); -- 
    req_1916_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1916_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(237), ack => WPIPE_Block0_start_974_inst_req_1); -- 
    -- CP-element group 238:  transition  input  output  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	237 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	239 
    -- CP-element group 238:  members (6) 
      -- CP-element group 238: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_974_update_completed_
      -- CP-element group 238: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_974_Update/$exit
      -- CP-element group 238: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_974_Update/ack
      -- CP-element group 238: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_977_sample_start_
      -- CP-element group 238: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_977_Sample/$entry
      -- CP-element group 238: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_977_Sample/req
      -- 
    ack_1917_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_974_inst_ack_1, ack => convTranspose_CP_39_elements(238)); -- 
    req_1925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(238), ack => WPIPE_Block0_start_977_inst_req_0); -- 
    -- CP-element group 239:  transition  input  output  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	238 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	240 
    -- CP-element group 239:  members (6) 
      -- CP-element group 239: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_977_sample_completed_
      -- CP-element group 239: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_977_update_start_
      -- CP-element group 239: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_977_Sample/$exit
      -- CP-element group 239: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_977_Sample/ack
      -- CP-element group 239: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_977_Update/$entry
      -- CP-element group 239: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_977_Update/req
      -- 
    ack_1926_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_977_inst_ack_0, ack => convTranspose_CP_39_elements(239)); -- 
    req_1930_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1930_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(239), ack => WPIPE_Block0_start_977_inst_req_1); -- 
    -- CP-element group 240:  transition  input  output  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	239 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	241 
    -- CP-element group 240:  members (6) 
      -- CP-element group 240: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_977_update_completed_
      -- CP-element group 240: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_977_Update/$exit
      -- CP-element group 240: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_977_Update/ack
      -- CP-element group 240: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_980_sample_start_
      -- CP-element group 240: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_980_Sample/$entry
      -- CP-element group 240: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_980_Sample/req
      -- 
    ack_1931_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_977_inst_ack_1, ack => convTranspose_CP_39_elements(240)); -- 
    req_1939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(240), ack => WPIPE_Block0_start_980_inst_req_0); -- 
    -- CP-element group 241:  transition  input  output  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	240 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	242 
    -- CP-element group 241:  members (6) 
      -- CP-element group 241: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_980_sample_completed_
      -- CP-element group 241: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_980_update_start_
      -- CP-element group 241: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_980_Sample/$exit
      -- CP-element group 241: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_980_Sample/ack
      -- CP-element group 241: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_980_Update/$entry
      -- CP-element group 241: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_980_Update/req
      -- 
    ack_1940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_980_inst_ack_0, ack => convTranspose_CP_39_elements(241)); -- 
    req_1944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(241), ack => WPIPE_Block0_start_980_inst_req_1); -- 
    -- CP-element group 242:  transition  input  output  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	241 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	243 
    -- CP-element group 242:  members (6) 
      -- CP-element group 242: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_980_update_completed_
      -- CP-element group 242: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_980_Update/$exit
      -- CP-element group 242: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_980_Update/ack
      -- CP-element group 242: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_983_sample_start_
      -- CP-element group 242: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_983_Sample/$entry
      -- CP-element group 242: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_983_Sample/req
      -- 
    ack_1945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_980_inst_ack_1, ack => convTranspose_CP_39_elements(242)); -- 
    req_1953_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1953_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(242), ack => WPIPE_Block0_start_983_inst_req_0); -- 
    -- CP-element group 243:  transition  input  output  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	242 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	244 
    -- CP-element group 243:  members (6) 
      -- CP-element group 243: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_983_sample_completed_
      -- CP-element group 243: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_983_update_start_
      -- CP-element group 243: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_983_Sample/$exit
      -- CP-element group 243: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_983_Sample/ack
      -- CP-element group 243: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_983_Update/$entry
      -- CP-element group 243: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_983_Update/req
      -- 
    ack_1954_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_983_inst_ack_0, ack => convTranspose_CP_39_elements(243)); -- 
    req_1958_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1958_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(243), ack => WPIPE_Block0_start_983_inst_req_1); -- 
    -- CP-element group 244:  transition  input  output  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	243 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	245 
    -- CP-element group 244:  members (6) 
      -- CP-element group 244: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_983_update_completed_
      -- CP-element group 244: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_983_Update/$exit
      -- CP-element group 244: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_983_Update/ack
      -- CP-element group 244: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_986_sample_start_
      -- CP-element group 244: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_986_Sample/$entry
      -- CP-element group 244: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_986_Sample/req
      -- 
    ack_1959_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_983_inst_ack_1, ack => convTranspose_CP_39_elements(244)); -- 
    req_1967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(244), ack => WPIPE_Block0_start_986_inst_req_0); -- 
    -- CP-element group 245:  transition  input  output  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	244 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	246 
    -- CP-element group 245:  members (6) 
      -- CP-element group 245: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_986_sample_completed_
      -- CP-element group 245: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_986_update_start_
      -- CP-element group 245: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_986_Sample/$exit
      -- CP-element group 245: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_986_Sample/ack
      -- CP-element group 245: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_986_Update/$entry
      -- CP-element group 245: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_986_Update/req
      -- 
    ack_1968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_986_inst_ack_0, ack => convTranspose_CP_39_elements(245)); -- 
    req_1972_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1972_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(245), ack => WPIPE_Block0_start_986_inst_req_1); -- 
    -- CP-element group 246:  transition  input  output  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	245 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	247 
    -- CP-element group 246:  members (6) 
      -- CP-element group 246: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_986_update_completed_
      -- CP-element group 246: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_986_Update/$exit
      -- CP-element group 246: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_986_Update/ack
      -- CP-element group 246: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_989_sample_start_
      -- CP-element group 246: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_989_Sample/$entry
      -- CP-element group 246: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_989_Sample/req
      -- 
    ack_1973_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_986_inst_ack_1, ack => convTranspose_CP_39_elements(246)); -- 
    req_1981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(246), ack => WPIPE_Block0_start_989_inst_req_0); -- 
    -- CP-element group 247:  transition  input  output  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	246 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	248 
    -- CP-element group 247:  members (6) 
      -- CP-element group 247: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_989_sample_completed_
      -- CP-element group 247: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_989_update_start_
      -- CP-element group 247: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_989_Sample/$exit
      -- CP-element group 247: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_989_Sample/ack
      -- CP-element group 247: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_989_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_989_Update/req
      -- 
    ack_1982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_989_inst_ack_0, ack => convTranspose_CP_39_elements(247)); -- 
    req_1986_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1986_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(247), ack => WPIPE_Block0_start_989_inst_req_1); -- 
    -- CP-element group 248:  transition  input  output  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	247 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	249 
    -- CP-element group 248:  members (6) 
      -- CP-element group 248: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_989_update_completed_
      -- CP-element group 248: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_989_Update/$exit
      -- CP-element group 248: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_989_Update/ack
      -- CP-element group 248: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_992_sample_start_
      -- CP-element group 248: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_992_Sample/$entry
      -- CP-element group 248: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_992_Sample/req
      -- 
    ack_1987_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_989_inst_ack_1, ack => convTranspose_CP_39_elements(248)); -- 
    req_1995_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1995_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(248), ack => WPIPE_Block0_start_992_inst_req_0); -- 
    -- CP-element group 249:  transition  input  output  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	248 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	250 
    -- CP-element group 249:  members (6) 
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_992_sample_completed_
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_992_update_start_
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_992_Sample/$exit
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_992_Sample/ack
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_992_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_992_Update/req
      -- 
    ack_1996_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_992_inst_ack_0, ack => convTranspose_CP_39_elements(249)); -- 
    req_2000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(249), ack => WPIPE_Block0_start_992_inst_req_1); -- 
    -- CP-element group 250:  transition  input  output  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	249 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	251 
    -- CP-element group 250:  members (6) 
      -- CP-element group 250: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_992_update_completed_
      -- CP-element group 250: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_992_Update/$exit
      -- CP-element group 250: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_992_Update/ack
      -- CP-element group 250: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_995_sample_start_
      -- CP-element group 250: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_995_Sample/$entry
      -- CP-element group 250: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_995_Sample/req
      -- 
    ack_2001_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_992_inst_ack_1, ack => convTranspose_CP_39_elements(250)); -- 
    req_2009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(250), ack => WPIPE_Block0_start_995_inst_req_0); -- 
    -- CP-element group 251:  transition  input  output  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	250 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	252 
    -- CP-element group 251:  members (6) 
      -- CP-element group 251: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_995_sample_completed_
      -- CP-element group 251: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_995_update_start_
      -- CP-element group 251: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_995_Sample/$exit
      -- CP-element group 251: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_995_Sample/ack
      -- CP-element group 251: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_995_Update/$entry
      -- CP-element group 251: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_995_Update/req
      -- 
    ack_2010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_995_inst_ack_0, ack => convTranspose_CP_39_elements(251)); -- 
    req_2014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(251), ack => WPIPE_Block0_start_995_inst_req_1); -- 
    -- CP-element group 252:  transition  input  output  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	251 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	253 
    -- CP-element group 252:  members (6) 
      -- CP-element group 252: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_995_update_completed_
      -- CP-element group 252: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_995_Update/$exit
      -- CP-element group 252: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_995_Update/ack
      -- CP-element group 252: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_998_sample_start_
      -- CP-element group 252: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_998_Sample/$entry
      -- CP-element group 252: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_998_Sample/req
      -- 
    ack_2015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_995_inst_ack_1, ack => convTranspose_CP_39_elements(252)); -- 
    req_2023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(252), ack => WPIPE_Block0_start_998_inst_req_0); -- 
    -- CP-element group 253:  transition  input  output  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	252 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	254 
    -- CP-element group 253:  members (6) 
      -- CP-element group 253: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_998_sample_completed_
      -- CP-element group 253: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_998_update_start_
      -- CP-element group 253: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_998_Sample/$exit
      -- CP-element group 253: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_998_Sample/ack
      -- CP-element group 253: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_998_Update/$entry
      -- CP-element group 253: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_998_Update/req
      -- 
    ack_2024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_998_inst_ack_0, ack => convTranspose_CP_39_elements(253)); -- 
    req_2028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(253), ack => WPIPE_Block0_start_998_inst_req_1); -- 
    -- CP-element group 254:  transition  input  output  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	253 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	255 
    -- CP-element group 254:  members (6) 
      -- CP-element group 254: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_998_update_completed_
      -- CP-element group 254: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_998_Update/$exit
      -- CP-element group 254: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_998_Update/ack
      -- CP-element group 254: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1002_sample_start_
      -- CP-element group 254: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1002_Sample/$entry
      -- CP-element group 254: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1002_Sample/req
      -- 
    ack_2029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_998_inst_ack_1, ack => convTranspose_CP_39_elements(254)); -- 
    req_2037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(254), ack => WPIPE_Block0_start_1002_inst_req_0); -- 
    -- CP-element group 255:  transition  input  output  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	254 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	256 
    -- CP-element group 255:  members (6) 
      -- CP-element group 255: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1002_Update/req
      -- CP-element group 255: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1002_Update/$entry
      -- CP-element group 255: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1002_sample_completed_
      -- CP-element group 255: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1002_update_start_
      -- CP-element group 255: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1002_Sample/$exit
      -- CP-element group 255: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1002_Sample/ack
      -- 
    ack_2038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1002_inst_ack_0, ack => convTranspose_CP_39_elements(255)); -- 
    req_2042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(255), ack => WPIPE_Block0_start_1002_inst_req_1); -- 
    -- CP-element group 256:  transition  input  output  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	255 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	257 
    -- CP-element group 256:  members (6) 
      -- CP-element group 256: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1006_sample_start_
      -- CP-element group 256: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1006_Sample/$entry
      -- CP-element group 256: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1006_Sample/req
      -- CP-element group 256: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1002_Update/ack
      -- CP-element group 256: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1002_Update/$exit
      -- CP-element group 256: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1002_update_completed_
      -- 
    ack_2043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1002_inst_ack_1, ack => convTranspose_CP_39_elements(256)); -- 
    req_2051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(256), ack => WPIPE_Block0_start_1006_inst_req_0); -- 
    -- CP-element group 257:  transition  input  output  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	256 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	258 
    -- CP-element group 257:  members (6) 
      -- CP-element group 257: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1006_Update/req
      -- CP-element group 257: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1006_Sample/$exit
      -- CP-element group 257: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1006_Sample/ack
      -- CP-element group 257: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1006_Update/$entry
      -- CP-element group 257: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1006_update_start_
      -- CP-element group 257: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1006_sample_completed_
      -- 
    ack_2052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1006_inst_ack_0, ack => convTranspose_CP_39_elements(257)); -- 
    req_2056_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2056_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(257), ack => WPIPE_Block0_start_1006_inst_req_1); -- 
    -- CP-element group 258:  transition  input  output  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	257 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	259 
    -- CP-element group 258:  members (6) 
      -- CP-element group 258: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1006_Update/$exit
      -- CP-element group 258: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1006_update_completed_
      -- CP-element group 258: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1006_Update/ack
      -- CP-element group 258: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1009_sample_start_
      -- CP-element group 258: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1009_Sample/$entry
      -- CP-element group 258: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1009_Sample/req
      -- 
    ack_2057_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1006_inst_ack_1, ack => convTranspose_CP_39_elements(258)); -- 
    req_2065_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2065_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(258), ack => WPIPE_Block0_start_1009_inst_req_0); -- 
    -- CP-element group 259:  transition  input  output  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	258 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	260 
    -- CP-element group 259:  members (6) 
      -- CP-element group 259: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1009_Update/req
      -- CP-element group 259: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1009_Sample/ack
      -- CP-element group 259: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1009_update_start_
      -- CP-element group 259: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1009_sample_completed_
      -- CP-element group 259: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1009_Sample/$exit
      -- CP-element group 259: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1009_Update/$entry
      -- 
    ack_2066_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1009_inst_ack_0, ack => convTranspose_CP_39_elements(259)); -- 
    req_2070_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2070_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(259), ack => WPIPE_Block0_start_1009_inst_req_1); -- 
    -- CP-element group 260:  transition  input  output  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	259 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	261 
    -- CP-element group 260:  members (6) 
      -- CP-element group 260: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1012_sample_start_
      -- CP-element group 260: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1012_Sample/$entry
      -- CP-element group 260: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1009_update_completed_
      -- CP-element group 260: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1009_Update/ack
      -- CP-element group 260: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1012_Sample/req
      -- CP-element group 260: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1009_Update/$exit
      -- 
    ack_2071_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1009_inst_ack_1, ack => convTranspose_CP_39_elements(260)); -- 
    req_2079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(260), ack => WPIPE_Block0_start_1012_inst_req_0); -- 
    -- CP-element group 261:  transition  input  output  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	260 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	262 
    -- CP-element group 261:  members (6) 
      -- CP-element group 261: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1012_sample_completed_
      -- CP-element group 261: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1012_Sample/$exit
      -- CP-element group 261: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1012_update_start_
      -- CP-element group 261: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1012_Sample/ack
      -- CP-element group 261: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1012_Update/$entry
      -- CP-element group 261: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1012_Update/req
      -- 
    ack_2080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1012_inst_ack_0, ack => convTranspose_CP_39_elements(261)); -- 
    req_2084_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2084_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(261), ack => WPIPE_Block0_start_1012_inst_req_1); -- 
    -- CP-element group 262:  transition  input  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	261 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	373 
    -- CP-element group 262:  members (3) 
      -- CP-element group 262: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1012_update_completed_
      -- CP-element group 262: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1012_Update/$exit
      -- CP-element group 262: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block0_start_1012_Update/ack
      -- 
    ack_2085_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1012_inst_ack_1, ack => convTranspose_CP_39_elements(262)); -- 
    -- CP-element group 263:  transition  input  output  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	234 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	264 
    -- CP-element group 263:  members (6) 
      -- CP-element group 263: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1015_Update/req
      -- CP-element group 263: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1015_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1015_Sample/ack
      -- CP-element group 263: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1015_Sample/$exit
      -- CP-element group 263: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1015_update_start_
      -- CP-element group 263: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1015_sample_completed_
      -- 
    ack_2094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1015_inst_ack_0, ack => convTranspose_CP_39_elements(263)); -- 
    req_2098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(263), ack => WPIPE_Block1_start_1015_inst_req_1); -- 
    -- CP-element group 264:  transition  input  output  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	263 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	265 
    -- CP-element group 264:  members (6) 
      -- CP-element group 264: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1018_Sample/req
      -- CP-element group 264: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1018_Sample/$entry
      -- CP-element group 264: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1018_sample_start_
      -- CP-element group 264: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1015_Update/ack
      -- CP-element group 264: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1015_Update/$exit
      -- CP-element group 264: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1015_update_completed_
      -- 
    ack_2099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1015_inst_ack_1, ack => convTranspose_CP_39_elements(264)); -- 
    req_2107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(264), ack => WPIPE_Block1_start_1018_inst_req_0); -- 
    -- CP-element group 265:  transition  input  output  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	264 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	266 
    -- CP-element group 265:  members (6) 
      -- CP-element group 265: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1018_Update/req
      -- CP-element group 265: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1018_Update/$entry
      -- CP-element group 265: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1018_Sample/ack
      -- CP-element group 265: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1018_Sample/$exit
      -- CP-element group 265: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1018_update_start_
      -- CP-element group 265: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1018_sample_completed_
      -- 
    ack_2108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1018_inst_ack_0, ack => convTranspose_CP_39_elements(265)); -- 
    req_2112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(265), ack => WPIPE_Block1_start_1018_inst_req_1); -- 
    -- CP-element group 266:  transition  input  output  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	265 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	267 
    -- CP-element group 266:  members (6) 
      -- CP-element group 266: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1018_Update/$exit
      -- CP-element group 266: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1018_Update/ack
      -- CP-element group 266: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1021_sample_start_
      -- CP-element group 266: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1021_Sample/req
      -- CP-element group 266: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1021_Sample/$entry
      -- CP-element group 266: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1018_update_completed_
      -- 
    ack_2113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1018_inst_ack_1, ack => convTranspose_CP_39_elements(266)); -- 
    req_2121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(266), ack => WPIPE_Block1_start_1021_inst_req_0); -- 
    -- CP-element group 267:  transition  input  output  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	266 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	268 
    -- CP-element group 267:  members (6) 
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1021_Sample/$exit
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1021_update_start_
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1021_sample_completed_
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1021_Sample/ack
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1021_Update/$entry
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1021_Update/req
      -- 
    ack_2122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1021_inst_ack_0, ack => convTranspose_CP_39_elements(267)); -- 
    req_2126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(267), ack => WPIPE_Block1_start_1021_inst_req_1); -- 
    -- CP-element group 268:  transition  input  output  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	267 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	269 
    -- CP-element group 268:  members (6) 
      -- CP-element group 268: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1021_update_completed_
      -- CP-element group 268: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1021_Update/ack
      -- CP-element group 268: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1024_sample_start_
      -- CP-element group 268: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1021_Update/$exit
      -- CP-element group 268: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1024_Sample/$entry
      -- CP-element group 268: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1024_Sample/req
      -- 
    ack_2127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1021_inst_ack_1, ack => convTranspose_CP_39_elements(268)); -- 
    req_2135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(268), ack => WPIPE_Block1_start_1024_inst_req_0); -- 
    -- CP-element group 269:  transition  input  output  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	268 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	270 
    -- CP-element group 269:  members (6) 
      -- CP-element group 269: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1024_sample_completed_
      -- CP-element group 269: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1024_update_start_
      -- CP-element group 269: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1024_Sample/$exit
      -- CP-element group 269: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1024_Sample/ack
      -- CP-element group 269: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1024_Update/$entry
      -- CP-element group 269: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1024_Update/req
      -- 
    ack_2136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 269_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1024_inst_ack_0, ack => convTranspose_CP_39_elements(269)); -- 
    req_2140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(269), ack => WPIPE_Block1_start_1024_inst_req_1); -- 
    -- CP-element group 270:  transition  input  output  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	269 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	271 
    -- CP-element group 270:  members (6) 
      -- CP-element group 270: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1024_update_completed_
      -- CP-element group 270: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1024_Update/$exit
      -- CP-element group 270: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1024_Update/ack
      -- CP-element group 270: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1027_sample_start_
      -- CP-element group 270: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1027_Sample/req
      -- CP-element group 270: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1027_Sample/$entry
      -- 
    ack_2141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1024_inst_ack_1, ack => convTranspose_CP_39_elements(270)); -- 
    req_2149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(270), ack => WPIPE_Block1_start_1027_inst_req_0); -- 
    -- CP-element group 271:  transition  input  output  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	270 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	272 
    -- CP-element group 271:  members (6) 
      -- CP-element group 271: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1027_Update/req
      -- CP-element group 271: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1027_Sample/ack
      -- CP-element group 271: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1027_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1027_sample_completed_
      -- CP-element group 271: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1027_update_start_
      -- CP-element group 271: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1027_Sample/$exit
      -- 
    ack_2150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1027_inst_ack_0, ack => convTranspose_CP_39_elements(271)); -- 
    req_2154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(271), ack => WPIPE_Block1_start_1027_inst_req_1); -- 
    -- CP-element group 272:  transition  input  output  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	271 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	273 
    -- CP-element group 272:  members (6) 
      -- CP-element group 272: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1027_Update/$exit
      -- CP-element group 272: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1027_Update/ack
      -- CP-element group 272: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1030_sample_start_
      -- CP-element group 272: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1027_update_completed_
      -- CP-element group 272: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1030_Sample/req
      -- CP-element group 272: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1030_Sample/$entry
      -- 
    ack_2155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1027_inst_ack_1, ack => convTranspose_CP_39_elements(272)); -- 
    req_2163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(272), ack => WPIPE_Block1_start_1030_inst_req_0); -- 
    -- CP-element group 273:  transition  input  output  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	272 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	274 
    -- CP-element group 273:  members (6) 
      -- CP-element group 273: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1030_sample_completed_
      -- CP-element group 273: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1030_Update/req
      -- CP-element group 273: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1030_Update/$entry
      -- CP-element group 273: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1030_Sample/ack
      -- CP-element group 273: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1030_Sample/$exit
      -- CP-element group 273: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1030_update_start_
      -- 
    ack_2164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1030_inst_ack_0, ack => convTranspose_CP_39_elements(273)); -- 
    req_2168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(273), ack => WPIPE_Block1_start_1030_inst_req_1); -- 
    -- CP-element group 274:  transition  input  output  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	273 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	275 
    -- CP-element group 274:  members (6) 
      -- CP-element group 274: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1033_Sample/req
      -- CP-element group 274: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1033_Sample/$entry
      -- CP-element group 274: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1033_sample_start_
      -- CP-element group 274: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1030_Update/ack
      -- CP-element group 274: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1030_Update/$exit
      -- CP-element group 274: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1030_update_completed_
      -- 
    ack_2169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1030_inst_ack_1, ack => convTranspose_CP_39_elements(274)); -- 
    req_2177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(274), ack => WPIPE_Block1_start_1033_inst_req_0); -- 
    -- CP-element group 275:  transition  input  output  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	274 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	276 
    -- CP-element group 275:  members (6) 
      -- CP-element group 275: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1033_Update/req
      -- CP-element group 275: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1033_Update/$entry
      -- CP-element group 275: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1033_Sample/ack
      -- CP-element group 275: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1033_Sample/$exit
      -- CP-element group 275: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1033_update_start_
      -- CP-element group 275: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1033_sample_completed_
      -- 
    ack_2178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1033_inst_ack_0, ack => convTranspose_CP_39_elements(275)); -- 
    req_2182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(275), ack => WPIPE_Block1_start_1033_inst_req_1); -- 
    -- CP-element group 276:  transition  input  output  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	275 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	277 
    -- CP-element group 276:  members (6) 
      -- CP-element group 276: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1036_Sample/req
      -- CP-element group 276: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1036_Sample/$entry
      -- CP-element group 276: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1036_sample_start_
      -- CP-element group 276: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1033_Update/ack
      -- CP-element group 276: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1033_Update/$exit
      -- CP-element group 276: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1033_update_completed_
      -- 
    ack_2183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1033_inst_ack_1, ack => convTranspose_CP_39_elements(276)); -- 
    req_2191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(276), ack => WPIPE_Block1_start_1036_inst_req_0); -- 
    -- CP-element group 277:  transition  input  output  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	276 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	278 
    -- CP-element group 277:  members (6) 
      -- CP-element group 277: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1036_Update/req
      -- CP-element group 277: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1036_Update/$entry
      -- CP-element group 277: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1036_Sample/ack
      -- CP-element group 277: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1036_Sample/$exit
      -- CP-element group 277: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1036_update_start_
      -- CP-element group 277: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1036_sample_completed_
      -- 
    ack_2192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1036_inst_ack_0, ack => convTranspose_CP_39_elements(277)); -- 
    req_2196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(277), ack => WPIPE_Block1_start_1036_inst_req_1); -- 
    -- CP-element group 278:  transition  input  output  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	277 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	279 
    -- CP-element group 278:  members (6) 
      -- CP-element group 278: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1039_Sample/req
      -- CP-element group 278: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1039_Sample/$entry
      -- CP-element group 278: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1039_sample_start_
      -- CP-element group 278: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1036_Update/ack
      -- CP-element group 278: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1036_Update/$exit
      -- CP-element group 278: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1036_update_completed_
      -- 
    ack_2197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1036_inst_ack_1, ack => convTranspose_CP_39_elements(278)); -- 
    req_2205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(278), ack => WPIPE_Block1_start_1039_inst_req_0); -- 
    -- CP-element group 279:  transition  input  output  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	278 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	280 
    -- CP-element group 279:  members (6) 
      -- CP-element group 279: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1039_Update/req
      -- CP-element group 279: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1039_Update/$entry
      -- CP-element group 279: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1039_Sample/ack
      -- CP-element group 279: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1039_Sample/$exit
      -- CP-element group 279: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1039_update_start_
      -- CP-element group 279: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1039_sample_completed_
      -- 
    ack_2206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1039_inst_ack_0, ack => convTranspose_CP_39_elements(279)); -- 
    req_2210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(279), ack => WPIPE_Block1_start_1039_inst_req_1); -- 
    -- CP-element group 280:  transition  input  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	279 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	283 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1039_Update/ack
      -- CP-element group 280: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1039_Update/$exit
      -- CP-element group 280: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1039_update_completed_
      -- 
    ack_2211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1039_inst_ack_1, ack => convTranspose_CP_39_elements(280)); -- 
    -- CP-element group 281:  transition  input  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	234 
    -- CP-element group 281: successors 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1050_Sample/ra
      -- CP-element group 281: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1050_sample_completed_
      -- CP-element group 281: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1050_Sample/$exit
      -- 
    ra_2220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1050_inst_ack_0, ack => convTranspose_CP_39_elements(281)); -- 
    -- CP-element group 282:  transition  input  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	234 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	283 
    -- CP-element group 282:  members (3) 
      -- CP-element group 282: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1050_Update/$exit
      -- CP-element group 282: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1050_update_completed_
      -- CP-element group 282: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1050_Update/ca
      -- 
    ca_2225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1050_inst_ack_1, ack => convTranspose_CP_39_elements(282)); -- 
    -- CP-element group 283:  join  transition  output  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	280 
    -- CP-element group 283: 	282 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	284 
    -- CP-element group 283:  members (3) 
      -- CP-element group 283: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1052_Sample/req
      -- CP-element group 283: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1052_sample_start_
      -- CP-element group 283: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1052_Sample/$entry
      -- 
    req_2233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(283), ack => WPIPE_Block1_start_1052_inst_req_0); -- 
    convTranspose_cp_element_group_283: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_283"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(280) & convTranspose_CP_39_elements(282);
      gj_convTranspose_cp_element_group_283 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(283), clk => clk, reset => reset); --
    end block;
    -- CP-element group 284:  transition  input  output  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	283 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	285 
    -- CP-element group 284:  members (6) 
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1052_Sample/ack
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1052_sample_completed_
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1052_update_start_
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1052_Sample/$exit
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1052_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1052_Update/req
      -- 
    ack_2234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1052_inst_ack_0, ack => convTranspose_CP_39_elements(284)); -- 
    req_2238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(284), ack => WPIPE_Block1_start_1052_inst_req_1); -- 
    -- CP-element group 285:  transition  input  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	284 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	288 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1052_update_completed_
      -- CP-element group 285: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1052_Update/$exit
      -- CP-element group 285: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1052_Update/ack
      -- 
    ack_2239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1052_inst_ack_1, ack => convTranspose_CP_39_elements(285)); -- 
    -- CP-element group 286:  transition  input  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	234 
    -- CP-element group 286: successors 
    -- CP-element group 286:  members (3) 
      -- CP-element group 286: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1057_sample_completed_
      -- CP-element group 286: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1057_Sample/$exit
      -- CP-element group 286: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1057_Sample/ra
      -- 
    ra_2248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1057_inst_ack_0, ack => convTranspose_CP_39_elements(286)); -- 
    -- CP-element group 287:  transition  input  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	234 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	288 
    -- CP-element group 287:  members (3) 
      -- CP-element group 287: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1057_update_completed_
      -- CP-element group 287: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1057_Update/ca
      -- CP-element group 287: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1057_Update/$exit
      -- 
    ca_2253_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1057_inst_ack_1, ack => convTranspose_CP_39_elements(287)); -- 
    -- CP-element group 288:  join  transition  output  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	285 
    -- CP-element group 288: 	287 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	289 
    -- CP-element group 288:  members (3) 
      -- CP-element group 288: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1059_Sample/req
      -- CP-element group 288: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1059_Sample/$entry
      -- CP-element group 288: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1059_sample_start_
      -- 
    req_2261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(288), ack => WPIPE_Block1_start_1059_inst_req_0); -- 
    convTranspose_cp_element_group_288: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_288"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(285) & convTranspose_CP_39_elements(287);
      gj_convTranspose_cp_element_group_288 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(288), clk => clk, reset => reset); --
    end block;
    -- CP-element group 289:  transition  input  output  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	288 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	290 
    -- CP-element group 289:  members (6) 
      -- CP-element group 289: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1059_Sample/$exit
      -- CP-element group 289: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1059_Sample/ack
      -- CP-element group 289: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1059_Update/req
      -- CP-element group 289: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1059_Update/$entry
      -- CP-element group 289: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1059_update_start_
      -- CP-element group 289: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1059_sample_completed_
      -- 
    ack_2262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1059_inst_ack_0, ack => convTranspose_CP_39_elements(289)); -- 
    req_2266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(289), ack => WPIPE_Block1_start_1059_inst_req_1); -- 
    -- CP-element group 290:  transition  input  output  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	289 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	291 
    -- CP-element group 290:  members (6) 
      -- CP-element group 290: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1059_Update/$exit
      -- CP-element group 290: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1062_sample_start_
      -- CP-element group 290: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1059_Update/ack
      -- CP-element group 290: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1062_Sample/req
      -- CP-element group 290: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1062_Sample/$entry
      -- CP-element group 290: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1059_update_completed_
      -- 
    ack_2267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1059_inst_ack_1, ack => convTranspose_CP_39_elements(290)); -- 
    req_2275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(290), ack => WPIPE_Block1_start_1062_inst_req_0); -- 
    -- CP-element group 291:  transition  input  output  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	290 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	292 
    -- CP-element group 291:  members (6) 
      -- CP-element group 291: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1062_sample_completed_
      -- CP-element group 291: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1062_update_start_
      -- CP-element group 291: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1062_Sample/$exit
      -- CP-element group 291: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1062_Update/req
      -- CP-element group 291: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1062_Update/$entry
      -- CP-element group 291: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1062_Sample/ack
      -- 
    ack_2276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1062_inst_ack_0, ack => convTranspose_CP_39_elements(291)); -- 
    req_2280_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2280_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(291), ack => WPIPE_Block1_start_1062_inst_req_1); -- 
    -- CP-element group 292:  transition  input  output  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	291 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	293 
    -- CP-element group 292:  members (6) 
      -- CP-element group 292: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1062_update_completed_
      -- CP-element group 292: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1065_Sample/req
      -- CP-element group 292: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1065_Sample/$entry
      -- CP-element group 292: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1065_sample_start_
      -- CP-element group 292: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1062_Update/ack
      -- CP-element group 292: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1062_Update/$exit
      -- 
    ack_2281_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1062_inst_ack_1, ack => convTranspose_CP_39_elements(292)); -- 
    req_2289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(292), ack => WPIPE_Block1_start_1065_inst_req_0); -- 
    -- CP-element group 293:  transition  input  output  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	292 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	294 
    -- CP-element group 293:  members (6) 
      -- CP-element group 293: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1065_Update/req
      -- CP-element group 293: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1065_Update/$entry
      -- CP-element group 293: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1065_Sample/ack
      -- CP-element group 293: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1065_Sample/$exit
      -- CP-element group 293: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1065_update_start_
      -- CP-element group 293: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1065_sample_completed_
      -- 
    ack_2290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 293_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1065_inst_ack_0, ack => convTranspose_CP_39_elements(293)); -- 
    req_2294_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2294_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(293), ack => WPIPE_Block1_start_1065_inst_req_1); -- 
    -- CP-element group 294:  transition  input  output  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	293 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	295 
    -- CP-element group 294:  members (6) 
      -- CP-element group 294: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1068_Sample/req
      -- CP-element group 294: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1068_Sample/$entry
      -- CP-element group 294: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1068_sample_start_
      -- CP-element group 294: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1065_Update/ack
      -- CP-element group 294: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1065_Update/$exit
      -- CP-element group 294: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1065_update_completed_
      -- 
    ack_2295_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 294_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1065_inst_ack_1, ack => convTranspose_CP_39_elements(294)); -- 
    req_2303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(294), ack => WPIPE_Block1_start_1068_inst_req_0); -- 
    -- CP-element group 295:  transition  input  output  bypass 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	294 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	296 
    -- CP-element group 295:  members (6) 
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1068_Update/req
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1068_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1068_Sample/ack
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1068_Sample/$exit
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1068_update_start_
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1068_sample_completed_
      -- 
    ack_2304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1068_inst_ack_0, ack => convTranspose_CP_39_elements(295)); -- 
    req_2308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(295), ack => WPIPE_Block1_start_1068_inst_req_1); -- 
    -- CP-element group 296:  transition  input  bypass 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	295 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	373 
    -- CP-element group 296:  members (3) 
      -- CP-element group 296: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1068_Update/ack
      -- CP-element group 296: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1068_Update/$exit
      -- CP-element group 296: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block1_start_1068_update_completed_
      -- 
    ack_2309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1068_inst_ack_1, ack => convTranspose_CP_39_elements(296)); -- 
    -- CP-element group 297:  transition  input  output  bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	234 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	298 
    -- CP-element group 297:  members (6) 
      -- CP-element group 297: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1071_update_start_
      -- CP-element group 297: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1071_sample_completed_
      -- CP-element group 297: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1071_Sample/$exit
      -- CP-element group 297: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1071_Sample/ack
      -- CP-element group 297: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1071_Update/$entry
      -- CP-element group 297: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1071_Update/req
      -- 
    ack_2318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1071_inst_ack_0, ack => convTranspose_CP_39_elements(297)); -- 
    req_2322_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2322_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(297), ack => WPIPE_Block2_start_1071_inst_req_1); -- 
    -- CP-element group 298:  transition  input  output  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	297 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	299 
    -- CP-element group 298:  members (6) 
      -- CP-element group 298: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1071_Update/$exit
      -- CP-element group 298: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1071_Update/ack
      -- CP-element group 298: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1074_sample_start_
      -- CP-element group 298: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1074_Sample/$entry
      -- CP-element group 298: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1074_Sample/req
      -- CP-element group 298: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1071_update_completed_
      -- 
    ack_2323_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 298_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1071_inst_ack_1, ack => convTranspose_CP_39_elements(298)); -- 
    req_2331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(298), ack => WPIPE_Block2_start_1074_inst_req_0); -- 
    -- CP-element group 299:  transition  input  output  bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	298 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	300 
    -- CP-element group 299:  members (6) 
      -- CP-element group 299: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1074_sample_completed_
      -- CP-element group 299: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1074_update_start_
      -- CP-element group 299: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1074_Sample/$exit
      -- CP-element group 299: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1074_Sample/ack
      -- CP-element group 299: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1074_Update/$entry
      -- CP-element group 299: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1074_Update/req
      -- 
    ack_2332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1074_inst_ack_0, ack => convTranspose_CP_39_elements(299)); -- 
    req_2336_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2336_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(299), ack => WPIPE_Block2_start_1074_inst_req_1); -- 
    -- CP-element group 300:  transition  input  output  bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	299 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	301 
    -- CP-element group 300:  members (6) 
      -- CP-element group 300: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1074_update_completed_
      -- CP-element group 300: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1074_Update/$exit
      -- CP-element group 300: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1074_Update/ack
      -- CP-element group 300: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1077_sample_start_
      -- CP-element group 300: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1077_Sample/req
      -- CP-element group 300: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1077_Sample/$entry
      -- 
    ack_2337_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1074_inst_ack_1, ack => convTranspose_CP_39_elements(300)); -- 
    req_2345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(300), ack => WPIPE_Block2_start_1077_inst_req_0); -- 
    -- CP-element group 301:  transition  input  output  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	300 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	302 
    -- CP-element group 301:  members (6) 
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1077_sample_completed_
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1077_Update/req
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1077_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1077_Sample/ack
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1077_Sample/$exit
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1077_update_start_
      -- 
    ack_2346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 301_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1077_inst_ack_0, ack => convTranspose_CP_39_elements(301)); -- 
    req_2350_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2350_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(301), ack => WPIPE_Block2_start_1077_inst_req_1); -- 
    -- CP-element group 302:  transition  input  output  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	301 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	303 
    -- CP-element group 302:  members (6) 
      -- CP-element group 302: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1080_sample_start_
      -- CP-element group 302: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1080_Sample/$entry
      -- CP-element group 302: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1080_Sample/req
      -- CP-element group 302: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1077_Update/ack
      -- CP-element group 302: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1077_Update/$exit
      -- CP-element group 302: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1077_update_completed_
      -- 
    ack_2351_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 302_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1077_inst_ack_1, ack => convTranspose_CP_39_elements(302)); -- 
    req_2359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(302), ack => WPIPE_Block2_start_1080_inst_req_0); -- 
    -- CP-element group 303:  transition  input  output  bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	302 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	304 
    -- CP-element group 303:  members (6) 
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1080_update_start_
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1080_Sample/$exit
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1080_sample_completed_
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1080_Sample/ack
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1080_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1080_Update/req
      -- 
    ack_2360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1080_inst_ack_0, ack => convTranspose_CP_39_elements(303)); -- 
    req_2364_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2364_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(303), ack => WPIPE_Block2_start_1080_inst_req_1); -- 
    -- CP-element group 304:  transition  input  output  bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	303 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	305 
    -- CP-element group 304:  members (6) 
      -- CP-element group 304: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1083_sample_start_
      -- CP-element group 304: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1080_update_completed_
      -- CP-element group 304: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1083_Sample/$entry
      -- CP-element group 304: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1083_Sample/req
      -- CP-element group 304: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1080_Update/$exit
      -- CP-element group 304: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1080_Update/ack
      -- 
    ack_2365_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1080_inst_ack_1, ack => convTranspose_CP_39_elements(304)); -- 
    req_2373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(304), ack => WPIPE_Block2_start_1083_inst_req_0); -- 
    -- CP-element group 305:  transition  input  output  bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	304 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	306 
    -- CP-element group 305:  members (6) 
      -- CP-element group 305: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1083_update_start_
      -- CP-element group 305: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1083_sample_completed_
      -- CP-element group 305: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1083_Sample/$exit
      -- CP-element group 305: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1083_Sample/ack
      -- CP-element group 305: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1083_Update/$entry
      -- CP-element group 305: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1083_Update/req
      -- 
    ack_2374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 305_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1083_inst_ack_0, ack => convTranspose_CP_39_elements(305)); -- 
    req_2378_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2378_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(305), ack => WPIPE_Block2_start_1083_inst_req_1); -- 
    -- CP-element group 306:  transition  input  output  bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	305 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	307 
    -- CP-element group 306:  members (6) 
      -- CP-element group 306: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1083_update_completed_
      -- CP-element group 306: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1083_Update/$exit
      -- CP-element group 306: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1086_sample_start_
      -- CP-element group 306: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1083_Update/ack
      -- CP-element group 306: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1086_Sample/req
      -- CP-element group 306: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1086_Sample/$entry
      -- 
    ack_2379_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1083_inst_ack_1, ack => convTranspose_CP_39_elements(306)); -- 
    req_2387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(306), ack => WPIPE_Block2_start_1086_inst_req_0); -- 
    -- CP-element group 307:  transition  input  output  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	306 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	308 
    -- CP-element group 307:  members (6) 
      -- CP-element group 307: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1086_Update/req
      -- CP-element group 307: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1086_Update/$entry
      -- CP-element group 307: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1086_Sample/ack
      -- CP-element group 307: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1086_Sample/$exit
      -- CP-element group 307: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1086_update_start_
      -- CP-element group 307: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1086_sample_completed_
      -- 
    ack_2388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1086_inst_ack_0, ack => convTranspose_CP_39_elements(307)); -- 
    req_2392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(307), ack => WPIPE_Block2_start_1086_inst_req_1); -- 
    -- CP-element group 308:  transition  input  output  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	307 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	309 
    -- CP-element group 308:  members (6) 
      -- CP-element group 308: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1089_sample_start_
      -- CP-element group 308: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1086_Update/ack
      -- CP-element group 308: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1089_Sample/req
      -- CP-element group 308: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1086_Update/$exit
      -- CP-element group 308: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1089_Sample/$entry
      -- CP-element group 308: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1086_update_completed_
      -- 
    ack_2393_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1086_inst_ack_1, ack => convTranspose_CP_39_elements(308)); -- 
    req_2401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(308), ack => WPIPE_Block2_start_1089_inst_req_0); -- 
    -- CP-element group 309:  transition  input  output  bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	308 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	310 
    -- CP-element group 309:  members (6) 
      -- CP-element group 309: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1089_sample_completed_
      -- CP-element group 309: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1089_update_start_
      -- CP-element group 309: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1089_Update/req
      -- CP-element group 309: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1089_Update/$entry
      -- CP-element group 309: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1089_Sample/ack
      -- CP-element group 309: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1089_Sample/$exit
      -- 
    ack_2402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 309_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1089_inst_ack_0, ack => convTranspose_CP_39_elements(309)); -- 
    req_2406_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2406_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(309), ack => WPIPE_Block2_start_1089_inst_req_1); -- 
    -- CP-element group 310:  transition  input  output  bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	309 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	311 
    -- CP-element group 310:  members (6) 
      -- CP-element group 310: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1092_sample_start_
      -- CP-element group 310: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1092_Sample/$entry
      -- CP-element group 310: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1092_Sample/req
      -- CP-element group 310: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1089_Update/ack
      -- CP-element group 310: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1089_Update/$exit
      -- CP-element group 310: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1089_update_completed_
      -- 
    ack_2407_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 310_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1089_inst_ack_1, ack => convTranspose_CP_39_elements(310)); -- 
    req_2415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(310), ack => WPIPE_Block2_start_1092_inst_req_0); -- 
    -- CP-element group 311:  transition  input  output  bypass 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	310 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	312 
    -- CP-element group 311:  members (6) 
      -- CP-element group 311: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1092_sample_completed_
      -- CP-element group 311: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1092_update_start_
      -- CP-element group 311: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1092_Sample/$exit
      -- CP-element group 311: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1092_Update/req
      -- CP-element group 311: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1092_Update/$entry
      -- CP-element group 311: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1092_Sample/ack
      -- 
    ack_2416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1092_inst_ack_0, ack => convTranspose_CP_39_elements(311)); -- 
    req_2420_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2420_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(311), ack => WPIPE_Block2_start_1092_inst_req_1); -- 
    -- CP-element group 312:  transition  input  output  bypass 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	311 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	313 
    -- CP-element group 312:  members (6) 
      -- CP-element group 312: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1092_update_completed_
      -- CP-element group 312: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1092_Update/ack
      -- CP-element group 312: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1095_Sample/req
      -- CP-element group 312: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1095_Sample/$entry
      -- CP-element group 312: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1092_Update/$exit
      -- CP-element group 312: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1095_sample_start_
      -- 
    ack_2421_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1092_inst_ack_1, ack => convTranspose_CP_39_elements(312)); -- 
    req_2429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(312), ack => WPIPE_Block2_start_1095_inst_req_0); -- 
    -- CP-element group 313:  transition  input  output  bypass 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	312 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	314 
    -- CP-element group 313:  members (6) 
      -- CP-element group 313: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1095_Update/$entry
      -- CP-element group 313: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1095_Sample/ack
      -- CP-element group 313: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1095_Update/req
      -- CP-element group 313: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1095_update_start_
      -- CP-element group 313: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1095_Sample/$exit
      -- CP-element group 313: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1095_sample_completed_
      -- 
    ack_2430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1095_inst_ack_0, ack => convTranspose_CP_39_elements(313)); -- 
    req_2434_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2434_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(313), ack => WPIPE_Block2_start_1095_inst_req_1); -- 
    -- CP-element group 314:  transition  input  bypass 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	313 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	317 
    -- CP-element group 314:  members (3) 
      -- CP-element group 314: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1095_Update/ack
      -- CP-element group 314: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1095_Update/$exit
      -- CP-element group 314: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1095_update_completed_
      -- 
    ack_2435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1095_inst_ack_1, ack => convTranspose_CP_39_elements(314)); -- 
    -- CP-element group 315:  transition  input  bypass 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	234 
    -- CP-element group 315: successors 
    -- CP-element group 315:  members (3) 
      -- CP-element group 315: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1106_sample_completed_
      -- CP-element group 315: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1106_Sample/$exit
      -- CP-element group 315: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1106_Sample/ra
      -- 
    ra_2444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1106_inst_ack_0, ack => convTranspose_CP_39_elements(315)); -- 
    -- CP-element group 316:  transition  input  bypass 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	234 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	317 
    -- CP-element group 316:  members (3) 
      -- CP-element group 316: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1106_update_completed_
      -- CP-element group 316: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1106_Update/$exit
      -- CP-element group 316: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1106_Update/ca
      -- 
    ca_2449_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1106_inst_ack_1, ack => convTranspose_CP_39_elements(316)); -- 
    -- CP-element group 317:  join  transition  output  bypass 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	314 
    -- CP-element group 317: 	316 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	318 
    -- CP-element group 317:  members (3) 
      -- CP-element group 317: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1108_sample_start_
      -- CP-element group 317: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1108_Sample/$entry
      -- CP-element group 317: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1108_Sample/req
      -- 
    req_2457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(317), ack => WPIPE_Block2_start_1108_inst_req_0); -- 
    convTranspose_cp_element_group_317: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_317"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(314) & convTranspose_CP_39_elements(316);
      gj_convTranspose_cp_element_group_317 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(317), clk => clk, reset => reset); --
    end block;
    -- CP-element group 318:  transition  input  output  bypass 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	317 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	319 
    -- CP-element group 318:  members (6) 
      -- CP-element group 318: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1108_sample_completed_
      -- CP-element group 318: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1108_update_start_
      -- CP-element group 318: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1108_Sample/$exit
      -- CP-element group 318: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1108_Sample/ack
      -- CP-element group 318: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1108_Update/$entry
      -- CP-element group 318: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1108_Update/req
      -- 
    ack_2458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 318_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1108_inst_ack_0, ack => convTranspose_CP_39_elements(318)); -- 
    req_2462_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2462_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(318), ack => WPIPE_Block2_start_1108_inst_req_1); -- 
    -- CP-element group 319:  transition  input  bypass 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	318 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	322 
    -- CP-element group 319:  members (3) 
      -- CP-element group 319: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1108_update_completed_
      -- CP-element group 319: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1108_Update/$exit
      -- CP-element group 319: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1108_Update/ack
      -- 
    ack_2463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 319_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1108_inst_ack_1, ack => convTranspose_CP_39_elements(319)); -- 
    -- CP-element group 320:  transition  input  bypass 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	234 
    -- CP-element group 320: successors 
    -- CP-element group 320:  members (3) 
      -- CP-element group 320: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1113_sample_completed_
      -- CP-element group 320: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1113_Sample/$exit
      -- CP-element group 320: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1113_Sample/ra
      -- 
    ra_2472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 320_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1113_inst_ack_0, ack => convTranspose_CP_39_elements(320)); -- 
    -- CP-element group 321:  transition  input  bypass 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	234 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	322 
    -- CP-element group 321:  members (3) 
      -- CP-element group 321: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1113_update_completed_
      -- CP-element group 321: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1113_Update/$exit
      -- CP-element group 321: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1113_Update/ca
      -- 
    ca_2477_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1113_inst_ack_1, ack => convTranspose_CP_39_elements(321)); -- 
    -- CP-element group 322:  join  transition  output  bypass 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	319 
    -- CP-element group 322: 	321 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	323 
    -- CP-element group 322:  members (3) 
      -- CP-element group 322: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1115_sample_start_
      -- CP-element group 322: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1115_Sample/$entry
      -- CP-element group 322: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1115_Sample/req
      -- 
    req_2485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(322), ack => WPIPE_Block2_start_1115_inst_req_0); -- 
    convTranspose_cp_element_group_322: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_322"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(319) & convTranspose_CP_39_elements(321);
      gj_convTranspose_cp_element_group_322 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(322), clk => clk, reset => reset); --
    end block;
    -- CP-element group 323:  transition  input  output  bypass 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	322 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	324 
    -- CP-element group 323:  members (6) 
      -- CP-element group 323: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1115_Update/$entry
      -- CP-element group 323: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1115_sample_completed_
      -- CP-element group 323: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1115_update_start_
      -- CP-element group 323: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1115_Sample/$exit
      -- CP-element group 323: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1115_Sample/ack
      -- CP-element group 323: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1115_Update/req
      -- 
    ack_2486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 323_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1115_inst_ack_0, ack => convTranspose_CP_39_elements(323)); -- 
    req_2490_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2490_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(323), ack => WPIPE_Block2_start_1115_inst_req_1); -- 
    -- CP-element group 324:  transition  input  output  bypass 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	323 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	325 
    -- CP-element group 324:  members (6) 
      -- CP-element group 324: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1115_Update/$exit
      -- CP-element group 324: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1115_update_completed_
      -- CP-element group 324: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1115_Update/ack
      -- CP-element group 324: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1118_sample_start_
      -- CP-element group 324: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1118_Sample/$entry
      -- CP-element group 324: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1118_Sample/req
      -- 
    ack_2491_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 324_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1115_inst_ack_1, ack => convTranspose_CP_39_elements(324)); -- 
    req_2499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(324), ack => WPIPE_Block2_start_1118_inst_req_0); -- 
    -- CP-element group 325:  transition  input  output  bypass 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	324 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	326 
    -- CP-element group 325:  members (6) 
      -- CP-element group 325: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1118_sample_completed_
      -- CP-element group 325: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1118_update_start_
      -- CP-element group 325: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1118_Sample/$exit
      -- CP-element group 325: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1118_Sample/ack
      -- CP-element group 325: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1118_Update/$entry
      -- CP-element group 325: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1118_Update/req
      -- 
    ack_2500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 325_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1118_inst_ack_0, ack => convTranspose_CP_39_elements(325)); -- 
    req_2504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(325), ack => WPIPE_Block2_start_1118_inst_req_1); -- 
    -- CP-element group 326:  transition  input  output  bypass 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	325 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	327 
    -- CP-element group 326:  members (6) 
      -- CP-element group 326: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1118_update_completed_
      -- CP-element group 326: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1118_Update/$exit
      -- CP-element group 326: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1118_Update/ack
      -- CP-element group 326: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1121_sample_start_
      -- CP-element group 326: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1121_Sample/$entry
      -- CP-element group 326: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1121_Sample/req
      -- 
    ack_2505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 326_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1118_inst_ack_1, ack => convTranspose_CP_39_elements(326)); -- 
    req_2513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(326), ack => WPIPE_Block2_start_1121_inst_req_0); -- 
    -- CP-element group 327:  transition  input  output  bypass 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	326 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	328 
    -- CP-element group 327:  members (6) 
      -- CP-element group 327: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1121_sample_completed_
      -- CP-element group 327: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1121_update_start_
      -- CP-element group 327: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1121_Sample/$exit
      -- CP-element group 327: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1121_Sample/ack
      -- CP-element group 327: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1121_Update/$entry
      -- CP-element group 327: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1121_Update/req
      -- 
    ack_2514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 327_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1121_inst_ack_0, ack => convTranspose_CP_39_elements(327)); -- 
    req_2518_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2518_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(327), ack => WPIPE_Block2_start_1121_inst_req_1); -- 
    -- CP-element group 328:  transition  input  output  bypass 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	327 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	329 
    -- CP-element group 328:  members (6) 
      -- CP-element group 328: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1121_update_completed_
      -- CP-element group 328: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1121_Update/$exit
      -- CP-element group 328: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1121_Update/ack
      -- CP-element group 328: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1124_sample_start_
      -- CP-element group 328: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1124_Sample/$entry
      -- CP-element group 328: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1124_Sample/req
      -- 
    ack_2519_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 328_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1121_inst_ack_1, ack => convTranspose_CP_39_elements(328)); -- 
    req_2527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(328), ack => WPIPE_Block2_start_1124_inst_req_0); -- 
    -- CP-element group 329:  transition  input  output  bypass 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	328 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	330 
    -- CP-element group 329:  members (6) 
      -- CP-element group 329: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1124_sample_completed_
      -- CP-element group 329: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1124_update_start_
      -- CP-element group 329: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1124_Sample/$exit
      -- CP-element group 329: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1124_Sample/ack
      -- CP-element group 329: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1124_Update/$entry
      -- CP-element group 329: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1124_Update/req
      -- 
    ack_2528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 329_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1124_inst_ack_0, ack => convTranspose_CP_39_elements(329)); -- 
    req_2532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(329), ack => WPIPE_Block2_start_1124_inst_req_1); -- 
    -- CP-element group 330:  transition  input  bypass 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	329 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	373 
    -- CP-element group 330:  members (3) 
      -- CP-element group 330: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1124_update_completed_
      -- CP-element group 330: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1124_Update/$exit
      -- CP-element group 330: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block2_start_1124_Update/ack
      -- 
    ack_2533_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 330_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1124_inst_ack_1, ack => convTranspose_CP_39_elements(330)); -- 
    -- CP-element group 331:  transition  input  output  bypass 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	234 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	332 
    -- CP-element group 331:  members (6) 
      -- CP-element group 331: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1127_sample_completed_
      -- CP-element group 331: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1127_update_start_
      -- CP-element group 331: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1127_Sample/$exit
      -- CP-element group 331: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1127_Sample/ack
      -- CP-element group 331: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1127_Update/$entry
      -- CP-element group 331: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1127_Update/req
      -- 
    ack_2542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 331_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1127_inst_ack_0, ack => convTranspose_CP_39_elements(331)); -- 
    req_2546_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2546_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(331), ack => WPIPE_Block3_start_1127_inst_req_1); -- 
    -- CP-element group 332:  transition  input  output  bypass 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	331 
    -- CP-element group 332: successors 
    -- CP-element group 332: 	333 
    -- CP-element group 332:  members (6) 
      -- CP-element group 332: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1127_update_completed_
      -- CP-element group 332: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1127_Update/$exit
      -- CP-element group 332: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1127_Update/ack
      -- CP-element group 332: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1130_sample_start_
      -- CP-element group 332: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1130_Sample/$entry
      -- CP-element group 332: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1130_Sample/req
      -- 
    ack_2547_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1127_inst_ack_1, ack => convTranspose_CP_39_elements(332)); -- 
    req_2555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(332), ack => WPIPE_Block3_start_1130_inst_req_0); -- 
    -- CP-element group 333:  transition  input  output  bypass 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	332 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	334 
    -- CP-element group 333:  members (6) 
      -- CP-element group 333: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1130_sample_completed_
      -- CP-element group 333: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1130_update_start_
      -- CP-element group 333: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1130_Sample/$exit
      -- CP-element group 333: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1130_Sample/ack
      -- CP-element group 333: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1130_Update/$entry
      -- CP-element group 333: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1130_Update/req
      -- 
    ack_2556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 333_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1130_inst_ack_0, ack => convTranspose_CP_39_elements(333)); -- 
    req_2560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(333), ack => WPIPE_Block3_start_1130_inst_req_1); -- 
    -- CP-element group 334:  transition  input  output  bypass 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	333 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	335 
    -- CP-element group 334:  members (6) 
      -- CP-element group 334: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1130_update_completed_
      -- CP-element group 334: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1130_Update/$exit
      -- CP-element group 334: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1130_Update/ack
      -- CP-element group 334: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1133_sample_start_
      -- CP-element group 334: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1133_Sample/$entry
      -- CP-element group 334: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1133_Sample/req
      -- 
    ack_2561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 334_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1130_inst_ack_1, ack => convTranspose_CP_39_elements(334)); -- 
    req_2569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(334), ack => WPIPE_Block3_start_1133_inst_req_0); -- 
    -- CP-element group 335:  transition  input  output  bypass 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	334 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	336 
    -- CP-element group 335:  members (6) 
      -- CP-element group 335: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1133_sample_completed_
      -- CP-element group 335: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1133_update_start_
      -- CP-element group 335: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1133_Sample/$exit
      -- CP-element group 335: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1133_Sample/ack
      -- CP-element group 335: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1133_Update/$entry
      -- CP-element group 335: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1133_Update/req
      -- 
    ack_2570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 335_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1133_inst_ack_0, ack => convTranspose_CP_39_elements(335)); -- 
    req_2574_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2574_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(335), ack => WPIPE_Block3_start_1133_inst_req_1); -- 
    -- CP-element group 336:  transition  input  output  bypass 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	335 
    -- CP-element group 336: successors 
    -- CP-element group 336: 	337 
    -- CP-element group 336:  members (6) 
      -- CP-element group 336: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1133_update_completed_
      -- CP-element group 336: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1133_Update/$exit
      -- CP-element group 336: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1133_Update/ack
      -- CP-element group 336: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1136_sample_start_
      -- CP-element group 336: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1136_Sample/$entry
      -- CP-element group 336: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1136_Sample/req
      -- 
    ack_2575_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1133_inst_ack_1, ack => convTranspose_CP_39_elements(336)); -- 
    req_2583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(336), ack => WPIPE_Block3_start_1136_inst_req_0); -- 
    -- CP-element group 337:  transition  input  output  bypass 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	336 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	338 
    -- CP-element group 337:  members (6) 
      -- CP-element group 337: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1136_sample_completed_
      -- CP-element group 337: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1136_update_start_
      -- CP-element group 337: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1136_Sample/$exit
      -- CP-element group 337: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1136_Sample/ack
      -- CP-element group 337: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1136_Update/$entry
      -- CP-element group 337: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1136_Update/req
      -- 
    ack_2584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1136_inst_ack_0, ack => convTranspose_CP_39_elements(337)); -- 
    req_2588_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2588_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(337), ack => WPIPE_Block3_start_1136_inst_req_1); -- 
    -- CP-element group 338:  transition  input  output  bypass 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	337 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	339 
    -- CP-element group 338:  members (6) 
      -- CP-element group 338: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1136_update_completed_
      -- CP-element group 338: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1136_Update/$exit
      -- CP-element group 338: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1136_Update/ack
      -- CP-element group 338: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1139_sample_start_
      -- CP-element group 338: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1139_Sample/$entry
      -- CP-element group 338: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1139_Sample/req
      -- 
    ack_2589_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 338_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1136_inst_ack_1, ack => convTranspose_CP_39_elements(338)); -- 
    req_2597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(338), ack => WPIPE_Block3_start_1139_inst_req_0); -- 
    -- CP-element group 339:  transition  input  output  bypass 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	338 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	340 
    -- CP-element group 339:  members (6) 
      -- CP-element group 339: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1139_sample_completed_
      -- CP-element group 339: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1139_update_start_
      -- CP-element group 339: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1139_Sample/$exit
      -- CP-element group 339: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1139_Sample/ack
      -- CP-element group 339: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1139_Update/$entry
      -- CP-element group 339: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1139_Update/req
      -- 
    ack_2598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 339_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1139_inst_ack_0, ack => convTranspose_CP_39_elements(339)); -- 
    req_2602_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2602_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(339), ack => WPIPE_Block3_start_1139_inst_req_1); -- 
    -- CP-element group 340:  transition  input  output  bypass 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	339 
    -- CP-element group 340: successors 
    -- CP-element group 340: 	341 
    -- CP-element group 340:  members (6) 
      -- CP-element group 340: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1139_update_completed_
      -- CP-element group 340: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1139_Update/$exit
      -- CP-element group 340: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1139_Update/ack
      -- CP-element group 340: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1142_sample_start_
      -- CP-element group 340: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1142_Sample/$entry
      -- CP-element group 340: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1142_Sample/req
      -- 
    ack_2603_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1139_inst_ack_1, ack => convTranspose_CP_39_elements(340)); -- 
    req_2611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(340), ack => WPIPE_Block3_start_1142_inst_req_0); -- 
    -- CP-element group 341:  transition  input  output  bypass 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	340 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	342 
    -- CP-element group 341:  members (6) 
      -- CP-element group 341: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1142_sample_completed_
      -- CP-element group 341: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1142_update_start_
      -- CP-element group 341: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1142_Sample/$exit
      -- CP-element group 341: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1142_Sample/ack
      -- CP-element group 341: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1142_Update/$entry
      -- CP-element group 341: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1142_Update/req
      -- 
    ack_2612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1142_inst_ack_0, ack => convTranspose_CP_39_elements(341)); -- 
    req_2616_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2616_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(341), ack => WPIPE_Block3_start_1142_inst_req_1); -- 
    -- CP-element group 342:  transition  input  output  bypass 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	341 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	343 
    -- CP-element group 342:  members (6) 
      -- CP-element group 342: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1142_update_completed_
      -- CP-element group 342: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1142_Update/$exit
      -- CP-element group 342: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1142_Update/ack
      -- CP-element group 342: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1145_sample_start_
      -- CP-element group 342: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1145_Sample/$entry
      -- CP-element group 342: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1145_Sample/req
      -- 
    ack_2617_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 342_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1142_inst_ack_1, ack => convTranspose_CP_39_elements(342)); -- 
    req_2625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(342), ack => WPIPE_Block3_start_1145_inst_req_0); -- 
    -- CP-element group 343:  transition  input  output  bypass 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	342 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	344 
    -- CP-element group 343:  members (6) 
      -- CP-element group 343: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1145_sample_completed_
      -- CP-element group 343: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1145_update_start_
      -- CP-element group 343: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1145_Sample/$exit
      -- CP-element group 343: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1145_Sample/ack
      -- CP-element group 343: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1145_Update/$entry
      -- CP-element group 343: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1145_Update/req
      -- 
    ack_2626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 343_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1145_inst_ack_0, ack => convTranspose_CP_39_elements(343)); -- 
    req_2630_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2630_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(343), ack => WPIPE_Block3_start_1145_inst_req_1); -- 
    -- CP-element group 344:  transition  input  output  bypass 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	343 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	345 
    -- CP-element group 344:  members (6) 
      -- CP-element group 344: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1145_update_completed_
      -- CP-element group 344: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1145_Update/$exit
      -- CP-element group 344: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1145_Update/ack
      -- CP-element group 344: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1148_sample_start_
      -- CP-element group 344: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1148_Sample/$entry
      -- CP-element group 344: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1148_Sample/req
      -- 
    ack_2631_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 344_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1145_inst_ack_1, ack => convTranspose_CP_39_elements(344)); -- 
    req_2639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(344), ack => WPIPE_Block3_start_1148_inst_req_0); -- 
    -- CP-element group 345:  transition  input  output  bypass 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	344 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	346 
    -- CP-element group 345:  members (6) 
      -- CP-element group 345: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1148_sample_completed_
      -- CP-element group 345: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1148_update_start_
      -- CP-element group 345: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1148_Sample/$exit
      -- CP-element group 345: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1148_Sample/ack
      -- CP-element group 345: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1148_Update/$entry
      -- CP-element group 345: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1148_Update/req
      -- 
    ack_2640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 345_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1148_inst_ack_0, ack => convTranspose_CP_39_elements(345)); -- 
    req_2644_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2644_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(345), ack => WPIPE_Block3_start_1148_inst_req_1); -- 
    -- CP-element group 346:  transition  input  output  bypass 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	345 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	347 
    -- CP-element group 346:  members (6) 
      -- CP-element group 346: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1148_update_completed_
      -- CP-element group 346: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1148_Update/$exit
      -- CP-element group 346: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1148_Update/ack
      -- CP-element group 346: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1151_sample_start_
      -- CP-element group 346: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1151_Sample/$entry
      -- CP-element group 346: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1151_Sample/req
      -- 
    ack_2645_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 346_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1148_inst_ack_1, ack => convTranspose_CP_39_elements(346)); -- 
    req_2653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(346), ack => WPIPE_Block3_start_1151_inst_req_0); -- 
    -- CP-element group 347:  transition  input  output  bypass 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	346 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	348 
    -- CP-element group 347:  members (6) 
      -- CP-element group 347: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1151_sample_completed_
      -- CP-element group 347: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1151_update_start_
      -- CP-element group 347: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1151_Sample/$exit
      -- CP-element group 347: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1151_Sample/ack
      -- CP-element group 347: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1151_Update/$entry
      -- CP-element group 347: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1151_Update/req
      -- 
    ack_2654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 347_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1151_inst_ack_0, ack => convTranspose_CP_39_elements(347)); -- 
    req_2658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(347), ack => WPIPE_Block3_start_1151_inst_req_1); -- 
    -- CP-element group 348:  transition  input  bypass 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	347 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	351 
    -- CP-element group 348:  members (3) 
      -- CP-element group 348: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1151_update_completed_
      -- CP-element group 348: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1151_Update/$exit
      -- CP-element group 348: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1151_Update/ack
      -- 
    ack_2659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 348_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1151_inst_ack_1, ack => convTranspose_CP_39_elements(348)); -- 
    -- CP-element group 349:  transition  input  bypass 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	234 
    -- CP-element group 349: successors 
    -- CP-element group 349:  members (3) 
      -- CP-element group 349: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1162_sample_completed_
      -- CP-element group 349: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1162_Sample/$exit
      -- CP-element group 349: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1162_Sample/ra
      -- 
    ra_2668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 349_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1162_inst_ack_0, ack => convTranspose_CP_39_elements(349)); -- 
    -- CP-element group 350:  transition  input  bypass 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	234 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	351 
    -- CP-element group 350:  members (3) 
      -- CP-element group 350: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1162_update_completed_
      -- CP-element group 350: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1162_Update/$exit
      -- CP-element group 350: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1162_Update/ca
      -- 
    ca_2673_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 350_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1162_inst_ack_1, ack => convTranspose_CP_39_elements(350)); -- 
    -- CP-element group 351:  join  transition  output  bypass 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	348 
    -- CP-element group 351: 	350 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	352 
    -- CP-element group 351:  members (3) 
      -- CP-element group 351: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1164_sample_start_
      -- CP-element group 351: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1164_Sample/$entry
      -- CP-element group 351: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1164_Sample/req
      -- 
    req_2681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(351), ack => WPIPE_Block3_start_1164_inst_req_0); -- 
    convTranspose_cp_element_group_351: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_351"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(348) & convTranspose_CP_39_elements(350);
      gj_convTranspose_cp_element_group_351 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(351), clk => clk, reset => reset); --
    end block;
    -- CP-element group 352:  transition  input  output  bypass 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	351 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	353 
    -- CP-element group 352:  members (6) 
      -- CP-element group 352: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1164_sample_completed_
      -- CP-element group 352: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1164_update_start_
      -- CP-element group 352: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1164_Sample/$exit
      -- CP-element group 352: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1164_Sample/ack
      -- CP-element group 352: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1164_Update/$entry
      -- CP-element group 352: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1164_Update/req
      -- 
    ack_2682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1164_inst_ack_0, ack => convTranspose_CP_39_elements(352)); -- 
    req_2686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(352), ack => WPIPE_Block3_start_1164_inst_req_1); -- 
    -- CP-element group 353:  transition  input  bypass 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	352 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	356 
    -- CP-element group 353:  members (3) 
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1164_update_completed_
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1164_Update/$exit
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1164_Update/ack
      -- 
    ack_2687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 353_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1164_inst_ack_1, ack => convTranspose_CP_39_elements(353)); -- 
    -- CP-element group 354:  transition  input  bypass 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	234 
    -- CP-element group 354: successors 
    -- CP-element group 354:  members (3) 
      -- CP-element group 354: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1169_sample_completed_
      -- CP-element group 354: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1169_Sample/$exit
      -- CP-element group 354: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1169_Sample/ra
      -- 
    ra_2696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 354_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1169_inst_ack_0, ack => convTranspose_CP_39_elements(354)); -- 
    -- CP-element group 355:  transition  input  bypass 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	234 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	356 
    -- CP-element group 355:  members (3) 
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1169_update_completed_
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1169_Update/$exit
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/type_cast_1169_Update/ca
      -- 
    ca_2701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 355_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1169_inst_ack_1, ack => convTranspose_CP_39_elements(355)); -- 
    -- CP-element group 356:  join  transition  output  bypass 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	353 
    -- CP-element group 356: 	355 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	357 
    -- CP-element group 356:  members (3) 
      -- CP-element group 356: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1171_sample_start_
      -- CP-element group 356: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1171_Sample/$entry
      -- CP-element group 356: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1171_Sample/req
      -- 
    req_2709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(356), ack => WPIPE_Block3_start_1171_inst_req_0); -- 
    convTranspose_cp_element_group_356: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_356"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(353) & convTranspose_CP_39_elements(355);
      gj_convTranspose_cp_element_group_356 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(356), clk => clk, reset => reset); --
    end block;
    -- CP-element group 357:  transition  input  output  bypass 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	356 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	358 
    -- CP-element group 357:  members (6) 
      -- CP-element group 357: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1171_sample_completed_
      -- CP-element group 357: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1171_update_start_
      -- CP-element group 357: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1171_Sample/$exit
      -- CP-element group 357: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1171_Sample/ack
      -- CP-element group 357: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1171_Update/$entry
      -- CP-element group 357: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1171_Update/req
      -- 
    ack_2710_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 357_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1171_inst_ack_0, ack => convTranspose_CP_39_elements(357)); -- 
    req_2714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(357), ack => WPIPE_Block3_start_1171_inst_req_1); -- 
    -- CP-element group 358:  transition  input  output  bypass 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	357 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	359 
    -- CP-element group 358:  members (6) 
      -- CP-element group 358: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1171_update_completed_
      -- CP-element group 358: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1171_Update/$exit
      -- CP-element group 358: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1171_Update/ack
      -- CP-element group 358: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1174_sample_start_
      -- CP-element group 358: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1174_Sample/$entry
      -- CP-element group 358: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1174_Sample/req
      -- 
    ack_2715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 358_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1171_inst_ack_1, ack => convTranspose_CP_39_elements(358)); -- 
    req_2723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(358), ack => WPIPE_Block3_start_1174_inst_req_0); -- 
    -- CP-element group 359:  transition  input  output  bypass 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	358 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	360 
    -- CP-element group 359:  members (6) 
      -- CP-element group 359: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1174_sample_completed_
      -- CP-element group 359: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1174_update_start_
      -- CP-element group 359: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1174_Sample/$exit
      -- CP-element group 359: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1174_Sample/ack
      -- CP-element group 359: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1174_Update/$entry
      -- CP-element group 359: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1174_Update/req
      -- 
    ack_2724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 359_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1174_inst_ack_0, ack => convTranspose_CP_39_elements(359)); -- 
    req_2728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(359), ack => WPIPE_Block3_start_1174_inst_req_1); -- 
    -- CP-element group 360:  transition  input  output  bypass 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	359 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	361 
    -- CP-element group 360:  members (6) 
      -- CP-element group 360: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1174_update_completed_
      -- CP-element group 360: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1174_Update/$exit
      -- CP-element group 360: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1174_Update/ack
      -- CP-element group 360: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1177_sample_start_
      -- CP-element group 360: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1177_Sample/$entry
      -- CP-element group 360: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1177_Sample/req
      -- 
    ack_2729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 360_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1174_inst_ack_1, ack => convTranspose_CP_39_elements(360)); -- 
    req_2737_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2737_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(360), ack => WPIPE_Block3_start_1177_inst_req_0); -- 
    -- CP-element group 361:  transition  input  output  bypass 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	360 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	362 
    -- CP-element group 361:  members (6) 
      -- CP-element group 361: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1177_sample_completed_
      -- CP-element group 361: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1177_update_start_
      -- CP-element group 361: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1177_Sample/$exit
      -- CP-element group 361: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1177_Sample/ack
      -- CP-element group 361: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1177_Update/$entry
      -- CP-element group 361: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1177_Update/req
      -- 
    ack_2738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 361_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1177_inst_ack_0, ack => convTranspose_CP_39_elements(361)); -- 
    req_2742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(361), ack => WPIPE_Block3_start_1177_inst_req_1); -- 
    -- CP-element group 362:  transition  input  output  bypass 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	361 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	363 
    -- CP-element group 362:  members (6) 
      -- CP-element group 362: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1177_update_completed_
      -- CP-element group 362: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1177_Update/$exit
      -- CP-element group 362: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1177_Update/ack
      -- CP-element group 362: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1180_sample_start_
      -- CP-element group 362: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1180_Sample/$entry
      -- CP-element group 362: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1180_Sample/req
      -- 
    ack_2743_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 362_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1177_inst_ack_1, ack => convTranspose_CP_39_elements(362)); -- 
    req_2751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(362), ack => WPIPE_Block3_start_1180_inst_req_0); -- 
    -- CP-element group 363:  transition  input  output  bypass 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	362 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	364 
    -- CP-element group 363:  members (6) 
      -- CP-element group 363: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1180_sample_completed_
      -- CP-element group 363: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1180_update_start_
      -- CP-element group 363: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1180_Sample/$exit
      -- CP-element group 363: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1180_Sample/ack
      -- CP-element group 363: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1180_Update/$entry
      -- CP-element group 363: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1180_Update/req
      -- 
    ack_2752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 363_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1180_inst_ack_0, ack => convTranspose_CP_39_elements(363)); -- 
    req_2756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(363), ack => WPIPE_Block3_start_1180_inst_req_1); -- 
    -- CP-element group 364:  transition  input  bypass 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	363 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	373 
    -- CP-element group 364:  members (3) 
      -- CP-element group 364: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1180_update_completed_
      -- CP-element group 364: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1180_Update/$exit
      -- CP-element group 364: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/WPIPE_Block3_start_1180_Update/ack
      -- 
    ack_2757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 364_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1180_inst_ack_1, ack => convTranspose_CP_39_elements(364)); -- 
    -- CP-element group 365:  transition  input  output  bypass 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	234 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	366 
    -- CP-element group 365:  members (6) 
      -- CP-element group 365: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block0_done_1184_sample_completed_
      -- CP-element group 365: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block0_done_1184_update_start_
      -- CP-element group 365: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block0_done_1184_Sample/$exit
      -- CP-element group 365: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block0_done_1184_Sample/ra
      -- CP-element group 365: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block0_done_1184_Update/$entry
      -- CP-element group 365: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block0_done_1184_Update/cr
      -- 
    ra_2766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 365_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1184_inst_ack_0, ack => convTranspose_CP_39_elements(365)); -- 
    cr_2770_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2770_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(365), ack => RPIPE_Block0_done_1184_inst_req_1); -- 
    -- CP-element group 366:  transition  input  bypass 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	365 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	373 
    -- CP-element group 366:  members (3) 
      -- CP-element group 366: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block0_done_1184_update_completed_
      -- CP-element group 366: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block0_done_1184_Update/$exit
      -- CP-element group 366: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block0_done_1184_Update/ca
      -- 
    ca_2771_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 366_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1184_inst_ack_1, ack => convTranspose_CP_39_elements(366)); -- 
    -- CP-element group 367:  transition  input  output  bypass 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	234 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	368 
    -- CP-element group 367:  members (6) 
      -- CP-element group 367: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block1_done_1187_sample_completed_
      -- CP-element group 367: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block1_done_1187_update_start_
      -- CP-element group 367: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block1_done_1187_Sample/$exit
      -- CP-element group 367: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block1_done_1187_Sample/ra
      -- CP-element group 367: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block1_done_1187_Update/$entry
      -- CP-element group 367: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block1_done_1187_Update/cr
      -- 
    ra_2780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 367_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1187_inst_ack_0, ack => convTranspose_CP_39_elements(367)); -- 
    cr_2784_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2784_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(367), ack => RPIPE_Block1_done_1187_inst_req_1); -- 
    -- CP-element group 368:  transition  input  bypass 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	367 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	373 
    -- CP-element group 368:  members (3) 
      -- CP-element group 368: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block1_done_1187_update_completed_
      -- CP-element group 368: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block1_done_1187_Update/$exit
      -- CP-element group 368: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block1_done_1187_Update/ca
      -- 
    ca_2785_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 368_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1187_inst_ack_1, ack => convTranspose_CP_39_elements(368)); -- 
    -- CP-element group 369:  transition  input  output  bypass 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	234 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	370 
    -- CP-element group 369:  members (6) 
      -- CP-element group 369: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block2_done_1190_sample_completed_
      -- CP-element group 369: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block2_done_1190_update_start_
      -- CP-element group 369: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block2_done_1190_Sample/$exit
      -- CP-element group 369: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block2_done_1190_Sample/ra
      -- CP-element group 369: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block2_done_1190_Update/$entry
      -- CP-element group 369: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block2_done_1190_Update/cr
      -- 
    ra_2794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 369_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1190_inst_ack_0, ack => convTranspose_CP_39_elements(369)); -- 
    cr_2798_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2798_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(369), ack => RPIPE_Block2_done_1190_inst_req_1); -- 
    -- CP-element group 370:  transition  input  bypass 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	369 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	373 
    -- CP-element group 370:  members (3) 
      -- CP-element group 370: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block2_done_1190_update_completed_
      -- CP-element group 370: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block2_done_1190_Update/$exit
      -- CP-element group 370: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block2_done_1190_Update/ca
      -- 
    ca_2799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 370_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1190_inst_ack_1, ack => convTranspose_CP_39_elements(370)); -- 
    -- CP-element group 371:  transition  input  output  bypass 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	234 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	372 
    -- CP-element group 371:  members (6) 
      -- CP-element group 371: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block3_done_1193_sample_completed_
      -- CP-element group 371: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block3_done_1193_update_start_
      -- CP-element group 371: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block3_done_1193_Sample/$exit
      -- CP-element group 371: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block3_done_1193_Sample/ra
      -- CP-element group 371: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block3_done_1193_Update/$entry
      -- CP-element group 371: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block3_done_1193_Update/cr
      -- 
    ra_2808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 371_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1193_inst_ack_0, ack => convTranspose_CP_39_elements(371)); -- 
    cr_2812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(371), ack => RPIPE_Block3_done_1193_inst_req_1); -- 
    -- CP-element group 372:  transition  input  bypass 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	371 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	373 
    -- CP-element group 372:  members (3) 
      -- CP-element group 372: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block3_done_1193_update_completed_
      -- CP-element group 372: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block3_done_1193_Update/$exit
      -- CP-element group 372: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/RPIPE_Block3_done_1193_Update/ca
      -- 
    ca_2813_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 372_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1193_inst_ack_1, ack => convTranspose_CP_39_elements(372)); -- 
    -- CP-element group 373:  join  fork  transition  place  output  bypass 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	330 
    -- CP-element group 373: 	364 
    -- CP-element group 373: 	366 
    -- CP-element group 373: 	368 
    -- CP-element group 373: 	370 
    -- CP-element group 373: 	372 
    -- CP-element group 373: 	262 
    -- CP-element group 373: 	296 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	374 
    -- CP-element group 373: 	375 
    -- CP-element group 373: 	377 
    -- CP-element group 373: 	381 
    -- CP-element group 373: 	383 
    -- CP-element group 373: 	385 
    -- CP-element group 373: 	387 
    -- CP-element group 373: 	389 
    -- CP-element group 373: 	391 
    -- CP-element group 373: 	393 
    -- CP-element group 373: 	395 
    -- CP-element group 373:  members (37) 
      -- CP-element group 373: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194__exit__
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308__entry__
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1283_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1283_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_33/assign_stmt_973_to_assign_stmt_1194/$exit
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/$entry
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/call_stmt_1197_sample_start_
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/call_stmt_1197_update_start_
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/call_stmt_1197_Sample/$entry
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/call_stmt_1197_Sample/crr
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/call_stmt_1197_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/call_stmt_1197_Update/ccr
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1201_update_start_
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1201_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1201_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1213_update_start_
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1213_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1213_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1223_update_start_
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1223_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1223_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1233_update_start_
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1233_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1233_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1243_update_start_
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1243_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1243_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1253_update_start_
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1253_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1253_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1263_update_start_
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1263_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1263_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1273_update_start_
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1273_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1273_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1283_update_start_
      -- 
    cr_2969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => type_cast_1283_inst_req_1); -- 
    crr_2824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => call_stmt_1197_call_req_0); -- 
    ccr_2829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => call_stmt_1197_call_req_1); -- 
    cr_2843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => type_cast_1201_inst_req_1); -- 
    cr_2871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => type_cast_1213_inst_req_1); -- 
    cr_2885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => type_cast_1223_inst_req_1); -- 
    cr_2899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => type_cast_1233_inst_req_1); -- 
    cr_2913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => type_cast_1243_inst_req_1); -- 
    cr_2927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => type_cast_1253_inst_req_1); -- 
    cr_2941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => type_cast_1263_inst_req_1); -- 
    cr_2955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => type_cast_1273_inst_req_1); -- 
    convTranspose_cp_element_group_373: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_373"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(330) & convTranspose_CP_39_elements(364) & convTranspose_CP_39_elements(366) & convTranspose_CP_39_elements(368) & convTranspose_CP_39_elements(370) & convTranspose_CP_39_elements(372) & convTranspose_CP_39_elements(262) & convTranspose_CP_39_elements(296);
      gj_convTranspose_cp_element_group_373 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(373), clk => clk, reset => reset); --
    end block;
    -- CP-element group 374:  transition  input  bypass 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	373 
    -- CP-element group 374: successors 
    -- CP-element group 374:  members (3) 
      -- CP-element group 374: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/call_stmt_1197_sample_completed_
      -- CP-element group 374: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/call_stmt_1197_Sample/$exit
      -- CP-element group 374: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/call_stmt_1197_Sample/cra
      -- 
    cra_2825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 374_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1197_call_ack_0, ack => convTranspose_CP_39_elements(374)); -- 
    -- CP-element group 375:  transition  input  output  bypass 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	373 
    -- CP-element group 375: successors 
    -- CP-element group 375: 	376 
    -- CP-element group 375:  members (6) 
      -- CP-element group 375: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/call_stmt_1197_update_completed_
      -- CP-element group 375: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/call_stmt_1197_Update/$exit
      -- CP-element group 375: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/call_stmt_1197_Update/cca
      -- CP-element group 375: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1201_sample_start_
      -- CP-element group 375: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1201_Sample/$entry
      -- CP-element group 375: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1201_Sample/rr
      -- 
    cca_2830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 375_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1197_call_ack_1, ack => convTranspose_CP_39_elements(375)); -- 
    rr_2838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(375), ack => type_cast_1201_inst_req_0); -- 
    -- CP-element group 376:  transition  input  bypass 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	375 
    -- CP-element group 376: successors 
    -- CP-element group 376:  members (3) 
      -- CP-element group 376: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1201_sample_completed_
      -- CP-element group 376: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1201_Sample/$exit
      -- CP-element group 376: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1201_Sample/ra
      -- 
    ra_2839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 376_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1201_inst_ack_0, ack => convTranspose_CP_39_elements(376)); -- 
    -- CP-element group 377:  fork  transition  input  output  bypass 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	373 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	378 
    -- CP-element group 377: 	380 
    -- CP-element group 377: 	382 
    -- CP-element group 377: 	384 
    -- CP-element group 377: 	386 
    -- CP-element group 377: 	388 
    -- CP-element group 377: 	390 
    -- CP-element group 377: 	392 
    -- CP-element group 377: 	394 
    -- CP-element group 377:  members (30) 
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1201_update_completed_
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1201_Update/$exit
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1201_Update/ca
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_elapsed_time_pipe_1208_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_elapsed_time_pipe_1208_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_elapsed_time_pipe_1208_Sample/req
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1213_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1213_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1213_Sample/rr
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1223_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1223_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1223_Sample/rr
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1233_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1233_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1233_Sample/rr
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1243_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1243_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1243_Sample/rr
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1253_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1253_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1253_Sample/rr
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1263_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1263_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1263_Sample/rr
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1273_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1273_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1273_Sample/rr
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1283_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1283_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1283_Sample/rr
      -- 
    ca_2844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 377_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1201_inst_ack_1, ack => convTranspose_CP_39_elements(377)); -- 
    req_2852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(377), ack => WPIPE_elapsed_time_pipe_1208_inst_req_0); -- 
    rr_2866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(377), ack => type_cast_1213_inst_req_0); -- 
    rr_2880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(377), ack => type_cast_1223_inst_req_0); -- 
    rr_2894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(377), ack => type_cast_1233_inst_req_0); -- 
    rr_2908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(377), ack => type_cast_1243_inst_req_0); -- 
    rr_2922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(377), ack => type_cast_1253_inst_req_0); -- 
    rr_2936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(377), ack => type_cast_1263_inst_req_0); -- 
    rr_2950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(377), ack => type_cast_1273_inst_req_0); -- 
    rr_2964_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2964_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(377), ack => type_cast_1283_inst_req_0); -- 
    -- CP-element group 378:  transition  input  output  bypass 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	377 
    -- CP-element group 378: successors 
    -- CP-element group 378: 	379 
    -- CP-element group 378:  members (6) 
      -- CP-element group 378: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_elapsed_time_pipe_1208_sample_completed_
      -- CP-element group 378: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_elapsed_time_pipe_1208_update_start_
      -- CP-element group 378: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_elapsed_time_pipe_1208_Sample/$exit
      -- CP-element group 378: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_elapsed_time_pipe_1208_Sample/ack
      -- CP-element group 378: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_elapsed_time_pipe_1208_Update/$entry
      -- CP-element group 378: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_elapsed_time_pipe_1208_Update/req
      -- 
    ack_2853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 378_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1208_inst_ack_0, ack => convTranspose_CP_39_elements(378)); -- 
    req_2857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(378), ack => WPIPE_elapsed_time_pipe_1208_inst_req_1); -- 
    -- CP-element group 379:  transition  input  bypass 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	378 
    -- CP-element group 379: successors 
    -- CP-element group 379: 	419 
    -- CP-element group 379:  members (3) 
      -- CP-element group 379: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_elapsed_time_pipe_1208_update_completed_
      -- CP-element group 379: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_elapsed_time_pipe_1208_Update/$exit
      -- CP-element group 379: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_elapsed_time_pipe_1208_Update/ack
      -- 
    ack_2858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 379_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1208_inst_ack_1, ack => convTranspose_CP_39_elements(379)); -- 
    -- CP-element group 380:  transition  input  bypass 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	377 
    -- CP-element group 380: successors 
    -- CP-element group 380:  members (3) 
      -- CP-element group 380: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1213_sample_completed_
      -- CP-element group 380: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1213_Sample/$exit
      -- CP-element group 380: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1213_Sample/ra
      -- 
    ra_2867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 380_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1213_inst_ack_0, ack => convTranspose_CP_39_elements(380)); -- 
    -- CP-element group 381:  transition  input  bypass 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	373 
    -- CP-element group 381: successors 
    -- CP-element group 381: 	416 
    -- CP-element group 381:  members (3) 
      -- CP-element group 381: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1213_update_completed_
      -- CP-element group 381: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1213_Update/$exit
      -- CP-element group 381: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1213_Update/ca
      -- 
    ca_2872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 381_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1213_inst_ack_1, ack => convTranspose_CP_39_elements(381)); -- 
    -- CP-element group 382:  transition  input  bypass 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	377 
    -- CP-element group 382: successors 
    -- CP-element group 382:  members (3) 
      -- CP-element group 382: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1223_sample_completed_
      -- CP-element group 382: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1223_Sample/$exit
      -- CP-element group 382: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1223_Sample/ra
      -- 
    ra_2881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 382_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1223_inst_ack_0, ack => convTranspose_CP_39_elements(382)); -- 
    -- CP-element group 383:  transition  input  bypass 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	373 
    -- CP-element group 383: successors 
    -- CP-element group 383: 	413 
    -- CP-element group 383:  members (3) 
      -- CP-element group 383: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1223_update_completed_
      -- CP-element group 383: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1223_Update/$exit
      -- CP-element group 383: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1223_Update/ca
      -- 
    ca_2886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 383_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1223_inst_ack_1, ack => convTranspose_CP_39_elements(383)); -- 
    -- CP-element group 384:  transition  input  bypass 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	377 
    -- CP-element group 384: successors 
    -- CP-element group 384:  members (3) 
      -- CP-element group 384: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1233_sample_completed_
      -- CP-element group 384: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1233_Sample/$exit
      -- CP-element group 384: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1233_Sample/ra
      -- 
    ra_2895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 384_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1233_inst_ack_0, ack => convTranspose_CP_39_elements(384)); -- 
    -- CP-element group 385:  transition  input  bypass 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	373 
    -- CP-element group 385: successors 
    -- CP-element group 385: 	410 
    -- CP-element group 385:  members (3) 
      -- CP-element group 385: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1233_update_completed_
      -- CP-element group 385: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1233_Update/$exit
      -- CP-element group 385: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1233_Update/ca
      -- 
    ca_2900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 385_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1233_inst_ack_1, ack => convTranspose_CP_39_elements(385)); -- 
    -- CP-element group 386:  transition  input  bypass 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	377 
    -- CP-element group 386: successors 
    -- CP-element group 386:  members (3) 
      -- CP-element group 386: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1243_sample_completed_
      -- CP-element group 386: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1243_Sample/$exit
      -- CP-element group 386: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1243_Sample/ra
      -- 
    ra_2909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 386_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1243_inst_ack_0, ack => convTranspose_CP_39_elements(386)); -- 
    -- CP-element group 387:  transition  input  bypass 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	373 
    -- CP-element group 387: successors 
    -- CP-element group 387: 	407 
    -- CP-element group 387:  members (3) 
      -- CP-element group 387: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1243_update_completed_
      -- CP-element group 387: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1243_Update/$exit
      -- CP-element group 387: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1243_Update/ca
      -- 
    ca_2914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 387_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1243_inst_ack_1, ack => convTranspose_CP_39_elements(387)); -- 
    -- CP-element group 388:  transition  input  bypass 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: 	377 
    -- CP-element group 388: successors 
    -- CP-element group 388:  members (3) 
      -- CP-element group 388: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1253_sample_completed_
      -- CP-element group 388: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1253_Sample/$exit
      -- CP-element group 388: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1253_Sample/ra
      -- 
    ra_2923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 388_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1253_inst_ack_0, ack => convTranspose_CP_39_elements(388)); -- 
    -- CP-element group 389:  transition  input  bypass 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	373 
    -- CP-element group 389: successors 
    -- CP-element group 389: 	404 
    -- CP-element group 389:  members (3) 
      -- CP-element group 389: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1253_update_completed_
      -- CP-element group 389: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1253_Update/$exit
      -- CP-element group 389: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1253_Update/ca
      -- 
    ca_2928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 389_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1253_inst_ack_1, ack => convTranspose_CP_39_elements(389)); -- 
    -- CP-element group 390:  transition  input  bypass 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: 	377 
    -- CP-element group 390: successors 
    -- CP-element group 390:  members (3) 
      -- CP-element group 390: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1263_sample_completed_
      -- CP-element group 390: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1263_Sample/$exit
      -- CP-element group 390: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1263_Sample/ra
      -- 
    ra_2937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 390_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1263_inst_ack_0, ack => convTranspose_CP_39_elements(390)); -- 
    -- CP-element group 391:  transition  input  bypass 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: 	373 
    -- CP-element group 391: successors 
    -- CP-element group 391: 	401 
    -- CP-element group 391:  members (3) 
      -- CP-element group 391: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1263_update_completed_
      -- CP-element group 391: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1263_Update/$exit
      -- CP-element group 391: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1263_Update/ca
      -- 
    ca_2942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 391_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1263_inst_ack_1, ack => convTranspose_CP_39_elements(391)); -- 
    -- CP-element group 392:  transition  input  bypass 
    -- CP-element group 392: predecessors 
    -- CP-element group 392: 	377 
    -- CP-element group 392: successors 
    -- CP-element group 392:  members (3) 
      -- CP-element group 392: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1273_sample_completed_
      -- CP-element group 392: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1273_Sample/$exit
      -- CP-element group 392: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1273_Sample/ra
      -- 
    ra_2951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 392_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1273_inst_ack_0, ack => convTranspose_CP_39_elements(392)); -- 
    -- CP-element group 393:  transition  input  bypass 
    -- CP-element group 393: predecessors 
    -- CP-element group 393: 	373 
    -- CP-element group 393: successors 
    -- CP-element group 393: 	398 
    -- CP-element group 393:  members (3) 
      -- CP-element group 393: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1273_update_completed_
      -- CP-element group 393: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1273_Update/$exit
      -- CP-element group 393: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1273_Update/ca
      -- 
    ca_2956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 393_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1273_inst_ack_1, ack => convTranspose_CP_39_elements(393)); -- 
    -- CP-element group 394:  transition  input  bypass 
    -- CP-element group 394: predecessors 
    -- CP-element group 394: 	377 
    -- CP-element group 394: successors 
    -- CP-element group 394:  members (3) 
      -- CP-element group 394: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1283_Sample/ra
      -- CP-element group 394: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1283_sample_completed_
      -- CP-element group 394: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1283_Sample/$exit
      -- 
    ra_2965_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 394_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1283_inst_ack_0, ack => convTranspose_CP_39_elements(394)); -- 
    -- CP-element group 395:  transition  input  output  bypass 
    -- CP-element group 395: predecessors 
    -- CP-element group 395: 	373 
    -- CP-element group 395: successors 
    -- CP-element group 395: 	396 
    -- CP-element group 395:  members (6) 
      -- CP-element group 395: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1283_Update/$exit
      -- CP-element group 395: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1283_Update/ca
      -- CP-element group 395: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1285_sample_start_
      -- CP-element group 395: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1285_Sample/$entry
      -- CP-element group 395: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1285_Sample/req
      -- CP-element group 395: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/type_cast_1283_update_completed_
      -- 
    ca_2970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 395_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1283_inst_ack_1, ack => convTranspose_CP_39_elements(395)); -- 
    req_2978_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2978_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(395), ack => WPIPE_ConvTranspose_output_pipe_1285_inst_req_0); -- 
    -- CP-element group 396:  transition  input  output  bypass 
    -- CP-element group 396: predecessors 
    -- CP-element group 396: 	395 
    -- CP-element group 396: successors 
    -- CP-element group 396: 	397 
    -- CP-element group 396:  members (6) 
      -- CP-element group 396: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1285_sample_completed_
      -- CP-element group 396: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1285_update_start_
      -- CP-element group 396: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1285_Sample/$exit
      -- CP-element group 396: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1285_Sample/ack
      -- CP-element group 396: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1285_Update/$entry
      -- CP-element group 396: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1285_Update/req
      -- 
    ack_2979_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 396_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1285_inst_ack_0, ack => convTranspose_CP_39_elements(396)); -- 
    req_2983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(396), ack => WPIPE_ConvTranspose_output_pipe_1285_inst_req_1); -- 
    -- CP-element group 397:  transition  input  bypass 
    -- CP-element group 397: predecessors 
    -- CP-element group 397: 	396 
    -- CP-element group 397: successors 
    -- CP-element group 397: 	398 
    -- CP-element group 397:  members (3) 
      -- CP-element group 397: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1285_update_completed_
      -- CP-element group 397: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1285_Update/$exit
      -- CP-element group 397: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1285_Update/ack
      -- 
    ack_2984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 397_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1285_inst_ack_1, ack => convTranspose_CP_39_elements(397)); -- 
    -- CP-element group 398:  join  transition  output  bypass 
    -- CP-element group 398: predecessors 
    -- CP-element group 398: 	393 
    -- CP-element group 398: 	397 
    -- CP-element group 398: successors 
    -- CP-element group 398: 	399 
    -- CP-element group 398:  members (3) 
      -- CP-element group 398: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1288_sample_start_
      -- CP-element group 398: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1288_Sample/req
      -- CP-element group 398: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1288_Sample/$entry
      -- 
    req_2992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(398), ack => WPIPE_ConvTranspose_output_pipe_1288_inst_req_0); -- 
    convTranspose_cp_element_group_398: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_398"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(393) & convTranspose_CP_39_elements(397);
      gj_convTranspose_cp_element_group_398 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(398), clk => clk, reset => reset); --
    end block;
    -- CP-element group 399:  transition  input  output  bypass 
    -- CP-element group 399: predecessors 
    -- CP-element group 399: 	398 
    -- CP-element group 399: successors 
    -- CP-element group 399: 	400 
    -- CP-element group 399:  members (6) 
      -- CP-element group 399: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1288_Sample/ack
      -- CP-element group 399: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1288_Update/$entry
      -- CP-element group 399: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1288_Update/req
      -- CP-element group 399: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1288_sample_completed_
      -- CP-element group 399: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1288_update_start_
      -- CP-element group 399: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1288_Sample/$exit
      -- 
    ack_2993_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 399_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1288_inst_ack_0, ack => convTranspose_CP_39_elements(399)); -- 
    req_2997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(399), ack => WPIPE_ConvTranspose_output_pipe_1288_inst_req_1); -- 
    -- CP-element group 400:  transition  input  bypass 
    -- CP-element group 400: predecessors 
    -- CP-element group 400: 	399 
    -- CP-element group 400: successors 
    -- CP-element group 400: 	401 
    -- CP-element group 400:  members (3) 
      -- CP-element group 400: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1288_Update/$exit
      -- CP-element group 400: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1288_Update/ack
      -- CP-element group 400: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1288_update_completed_
      -- 
    ack_2998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 400_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1288_inst_ack_1, ack => convTranspose_CP_39_elements(400)); -- 
    -- CP-element group 401:  join  transition  output  bypass 
    -- CP-element group 401: predecessors 
    -- CP-element group 401: 	391 
    -- CP-element group 401: 	400 
    -- CP-element group 401: successors 
    -- CP-element group 401: 	402 
    -- CP-element group 401:  members (3) 
      -- CP-element group 401: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1291_sample_start_
      -- CP-element group 401: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1291_Sample/req
      -- CP-element group 401: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1291_Sample/$entry
      -- 
    req_3006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(401), ack => WPIPE_ConvTranspose_output_pipe_1291_inst_req_0); -- 
    convTranspose_cp_element_group_401: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_401"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(391) & convTranspose_CP_39_elements(400);
      gj_convTranspose_cp_element_group_401 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(401), clk => clk, reset => reset); --
    end block;
    -- CP-element group 402:  transition  input  output  bypass 
    -- CP-element group 402: predecessors 
    -- CP-element group 402: 	401 
    -- CP-element group 402: successors 
    -- CP-element group 402: 	403 
    -- CP-element group 402:  members (6) 
      -- CP-element group 402: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1291_sample_completed_
      -- CP-element group 402: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1291_Update/req
      -- CP-element group 402: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1291_Update/$entry
      -- CP-element group 402: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1291_Sample/ack
      -- CP-element group 402: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1291_Sample/$exit
      -- CP-element group 402: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1291_update_start_
      -- 
    ack_3007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 402_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1291_inst_ack_0, ack => convTranspose_CP_39_elements(402)); -- 
    req_3011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(402), ack => WPIPE_ConvTranspose_output_pipe_1291_inst_req_1); -- 
    -- CP-element group 403:  transition  input  bypass 
    -- CP-element group 403: predecessors 
    -- CP-element group 403: 	402 
    -- CP-element group 403: successors 
    -- CP-element group 403: 	404 
    -- CP-element group 403:  members (3) 
      -- CP-element group 403: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1291_Update/ack
      -- CP-element group 403: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1291_Update/$exit
      -- CP-element group 403: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1291_update_completed_
      -- 
    ack_3012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 403_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1291_inst_ack_1, ack => convTranspose_CP_39_elements(403)); -- 
    -- CP-element group 404:  join  transition  output  bypass 
    -- CP-element group 404: predecessors 
    -- CP-element group 404: 	389 
    -- CP-element group 404: 	403 
    -- CP-element group 404: successors 
    -- CP-element group 404: 	405 
    -- CP-element group 404:  members (3) 
      -- CP-element group 404: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1294_Sample/req
      -- CP-element group 404: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1294_Sample/$entry
      -- CP-element group 404: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1294_sample_start_
      -- 
    req_3020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => WPIPE_ConvTranspose_output_pipe_1294_inst_req_0); -- 
    convTranspose_cp_element_group_404: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_404"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(389) & convTranspose_CP_39_elements(403);
      gj_convTranspose_cp_element_group_404 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(404), clk => clk, reset => reset); --
    end block;
    -- CP-element group 405:  transition  input  output  bypass 
    -- CP-element group 405: predecessors 
    -- CP-element group 405: 	404 
    -- CP-element group 405: successors 
    -- CP-element group 405: 	406 
    -- CP-element group 405:  members (6) 
      -- CP-element group 405: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1294_Update/req
      -- CP-element group 405: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1294_Update/$entry
      -- CP-element group 405: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1294_Sample/ack
      -- CP-element group 405: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1294_Sample/$exit
      -- CP-element group 405: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1294_update_start_
      -- CP-element group 405: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1294_sample_completed_
      -- 
    ack_3021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 405_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1294_inst_ack_0, ack => convTranspose_CP_39_elements(405)); -- 
    req_3025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(405), ack => WPIPE_ConvTranspose_output_pipe_1294_inst_req_1); -- 
    -- CP-element group 406:  transition  input  bypass 
    -- CP-element group 406: predecessors 
    -- CP-element group 406: 	405 
    -- CP-element group 406: successors 
    -- CP-element group 406: 	407 
    -- CP-element group 406:  members (3) 
      -- CP-element group 406: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1294_Update/ack
      -- CP-element group 406: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1294_Update/$exit
      -- CP-element group 406: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1294_update_completed_
      -- 
    ack_3026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 406_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1294_inst_ack_1, ack => convTranspose_CP_39_elements(406)); -- 
    -- CP-element group 407:  join  transition  output  bypass 
    -- CP-element group 407: predecessors 
    -- CP-element group 407: 	387 
    -- CP-element group 407: 	406 
    -- CP-element group 407: successors 
    -- CP-element group 407: 	408 
    -- CP-element group 407:  members (3) 
      -- CP-element group 407: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1297_Sample/req
      -- CP-element group 407: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1297_Sample/$entry
      -- CP-element group 407: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1297_sample_start_
      -- 
    req_3034_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3034_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(407), ack => WPIPE_ConvTranspose_output_pipe_1297_inst_req_0); -- 
    convTranspose_cp_element_group_407: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_407"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(387) & convTranspose_CP_39_elements(406);
      gj_convTranspose_cp_element_group_407 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(407), clk => clk, reset => reset); --
    end block;
    -- CP-element group 408:  transition  input  output  bypass 
    -- CP-element group 408: predecessors 
    -- CP-element group 408: 	407 
    -- CP-element group 408: successors 
    -- CP-element group 408: 	409 
    -- CP-element group 408:  members (6) 
      -- CP-element group 408: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1297_Update/req
      -- CP-element group 408: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1297_Update/$entry
      -- CP-element group 408: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1297_Sample/ack
      -- CP-element group 408: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1297_Sample/$exit
      -- CP-element group 408: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1297_update_start_
      -- CP-element group 408: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1297_sample_completed_
      -- 
    ack_3035_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 408_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1297_inst_ack_0, ack => convTranspose_CP_39_elements(408)); -- 
    req_3039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(408), ack => WPIPE_ConvTranspose_output_pipe_1297_inst_req_1); -- 
    -- CP-element group 409:  transition  input  bypass 
    -- CP-element group 409: predecessors 
    -- CP-element group 409: 	408 
    -- CP-element group 409: successors 
    -- CP-element group 409: 	410 
    -- CP-element group 409:  members (3) 
      -- CP-element group 409: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1297_Update/ack
      -- CP-element group 409: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1297_Update/$exit
      -- CP-element group 409: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1297_update_completed_
      -- 
    ack_3040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 409_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1297_inst_ack_1, ack => convTranspose_CP_39_elements(409)); -- 
    -- CP-element group 410:  join  transition  output  bypass 
    -- CP-element group 410: predecessors 
    -- CP-element group 410: 	385 
    -- CP-element group 410: 	409 
    -- CP-element group 410: successors 
    -- CP-element group 410: 	411 
    -- CP-element group 410:  members (3) 
      -- CP-element group 410: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1300_Sample/$entry
      -- CP-element group 410: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1300_Sample/req
      -- CP-element group 410: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1300_sample_start_
      -- 
    req_3048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(410), ack => WPIPE_ConvTranspose_output_pipe_1300_inst_req_0); -- 
    convTranspose_cp_element_group_410: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_410"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(385) & convTranspose_CP_39_elements(409);
      gj_convTranspose_cp_element_group_410 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(410), clk => clk, reset => reset); --
    end block;
    -- CP-element group 411:  transition  input  output  bypass 
    -- CP-element group 411: predecessors 
    -- CP-element group 411: 	410 
    -- CP-element group 411: successors 
    -- CP-element group 411: 	412 
    -- CP-element group 411:  members (6) 
      -- CP-element group 411: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1300_update_start_
      -- CP-element group 411: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1300_Sample/$exit
      -- CP-element group 411: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1300_Sample/ack
      -- CP-element group 411: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1300_Update/$entry
      -- CP-element group 411: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1300_Update/req
      -- CP-element group 411: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1300_sample_completed_
      -- 
    ack_3049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 411_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1300_inst_ack_0, ack => convTranspose_CP_39_elements(411)); -- 
    req_3053_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3053_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(411), ack => WPIPE_ConvTranspose_output_pipe_1300_inst_req_1); -- 
    -- CP-element group 412:  transition  input  bypass 
    -- CP-element group 412: predecessors 
    -- CP-element group 412: 	411 
    -- CP-element group 412: successors 
    -- CP-element group 412: 	413 
    -- CP-element group 412:  members (3) 
      -- CP-element group 412: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1300_update_completed_
      -- CP-element group 412: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1300_Update/$exit
      -- CP-element group 412: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1300_Update/ack
      -- 
    ack_3054_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 412_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1300_inst_ack_1, ack => convTranspose_CP_39_elements(412)); -- 
    -- CP-element group 413:  join  transition  output  bypass 
    -- CP-element group 413: predecessors 
    -- CP-element group 413: 	383 
    -- CP-element group 413: 	412 
    -- CP-element group 413: successors 
    -- CP-element group 413: 	414 
    -- CP-element group 413:  members (3) 
      -- CP-element group 413: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1303_sample_start_
      -- CP-element group 413: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1303_Sample/$entry
      -- CP-element group 413: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1303_Sample/req
      -- 
    req_3062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(413), ack => WPIPE_ConvTranspose_output_pipe_1303_inst_req_0); -- 
    convTranspose_cp_element_group_413: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_413"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(383) & convTranspose_CP_39_elements(412);
      gj_convTranspose_cp_element_group_413 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(413), clk => clk, reset => reset); --
    end block;
    -- CP-element group 414:  transition  input  output  bypass 
    -- CP-element group 414: predecessors 
    -- CP-element group 414: 	413 
    -- CP-element group 414: successors 
    -- CP-element group 414: 	415 
    -- CP-element group 414:  members (6) 
      -- CP-element group 414: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1303_Update/req
      -- CP-element group 414: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1303_sample_completed_
      -- CP-element group 414: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1303_update_start_
      -- CP-element group 414: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1303_Sample/$exit
      -- CP-element group 414: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1303_Sample/ack
      -- CP-element group 414: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1303_Update/$entry
      -- 
    ack_3063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 414_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1303_inst_ack_0, ack => convTranspose_CP_39_elements(414)); -- 
    req_3067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(414), ack => WPIPE_ConvTranspose_output_pipe_1303_inst_req_1); -- 
    -- CP-element group 415:  transition  input  bypass 
    -- CP-element group 415: predecessors 
    -- CP-element group 415: 	414 
    -- CP-element group 415: successors 
    -- CP-element group 415: 	416 
    -- CP-element group 415:  members (3) 
      -- CP-element group 415: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1303_Update/ack
      -- CP-element group 415: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1303_update_completed_
      -- CP-element group 415: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1303_Update/$exit
      -- 
    ack_3068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 415_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1303_inst_ack_1, ack => convTranspose_CP_39_elements(415)); -- 
    -- CP-element group 416:  join  transition  output  bypass 
    -- CP-element group 416: predecessors 
    -- CP-element group 416: 	381 
    -- CP-element group 416: 	415 
    -- CP-element group 416: successors 
    -- CP-element group 416: 	417 
    -- CP-element group 416:  members (3) 
      -- CP-element group 416: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1306_sample_start_
      -- CP-element group 416: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1306_Sample/req
      -- CP-element group 416: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1306_Sample/$entry
      -- 
    req_3076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(416), ack => WPIPE_ConvTranspose_output_pipe_1306_inst_req_0); -- 
    convTranspose_cp_element_group_416: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_416"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(381) & convTranspose_CP_39_elements(415);
      gj_convTranspose_cp_element_group_416 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(416), clk => clk, reset => reset); --
    end block;
    -- CP-element group 417:  transition  input  output  bypass 
    -- CP-element group 417: predecessors 
    -- CP-element group 417: 	416 
    -- CP-element group 417: successors 
    -- CP-element group 417: 	418 
    -- CP-element group 417:  members (6) 
      -- CP-element group 417: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1306_Update/req
      -- CP-element group 417: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1306_Update/$entry
      -- CP-element group 417: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1306_Sample/ack
      -- CP-element group 417: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1306_Sample/$exit
      -- CP-element group 417: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1306_update_start_
      -- CP-element group 417: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1306_sample_completed_
      -- 
    ack_3077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 417_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1306_inst_ack_0, ack => convTranspose_CP_39_elements(417)); -- 
    req_3081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(417), ack => WPIPE_ConvTranspose_output_pipe_1306_inst_req_1); -- 
    -- CP-element group 418:  transition  input  bypass 
    -- CP-element group 418: predecessors 
    -- CP-element group 418: 	417 
    -- CP-element group 418: successors 
    -- CP-element group 418: 	419 
    -- CP-element group 418:  members (3) 
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1306_Update/ack
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1306_Update/$exit
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/WPIPE_ConvTranspose_output_pipe_1306_update_completed_
      -- 
    ack_3082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 418_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1306_inst_ack_1, ack => convTranspose_CP_39_elements(418)); -- 
    -- CP-element group 419:  branch  join  transition  place  output  bypass 
    -- CP-element group 419: predecessors 
    -- CP-element group 419: 	379 
    -- CP-element group 419: 	418 
    -- CP-element group 419: successors 
    -- CP-element group 419: 	420 
    -- CP-element group 419: 	421 
    -- CP-element group 419:  members (10) 
      -- CP-element group 419: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308__exit__
      -- CP-element group 419: 	 branch_block_stmt_33/if_stmt_1310__entry__
      -- CP-element group 419: 	 branch_block_stmt_33/if_stmt_1310_else_link/$entry
      -- CP-element group 419: 	 branch_block_stmt_33/if_stmt_1310_if_link/$entry
      -- CP-element group 419: 	 branch_block_stmt_33/if_stmt_1310_eval_test/branch_req
      -- CP-element group 419: 	 branch_block_stmt_33/if_stmt_1310_eval_test/$exit
      -- CP-element group 419: 	 branch_block_stmt_33/if_stmt_1310_eval_test/$entry
      -- CP-element group 419: 	 branch_block_stmt_33/if_stmt_1310_dead_link/$entry
      -- CP-element group 419: 	 branch_block_stmt_33/R_cmp264506_1311_place
      -- CP-element group 419: 	 branch_block_stmt_33/call_stmt_1197_to_assign_stmt_1308/$exit
      -- 
    branch_req_3090_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3090_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(419), ack => if_stmt_1310_branch_req_0); -- 
    convTranspose_cp_element_group_419: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_419"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(379) & convTranspose_CP_39_elements(418);
      gj_convTranspose_cp_element_group_419 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(419), clk => clk, reset => reset); --
    end block;
    -- CP-element group 420:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 420: predecessors 
    -- CP-element group 420: 	419 
    -- CP-element group 420: successors 
    -- CP-element group 420: 	422 
    -- CP-element group 420: 	423 
    -- CP-element group 420:  members (18) 
      -- CP-element group 420: 	 branch_block_stmt_33/merge_stmt_1316__exit__
      -- CP-element group 420: 	 branch_block_stmt_33/assign_stmt_1322_to_assign_stmt_1351__entry__
      -- CP-element group 420: 	 branch_block_stmt_33/assign_stmt_1322_to_assign_stmt_1351/type_cast_1337_Update/cr
      -- CP-element group 420: 	 branch_block_stmt_33/assign_stmt_1322_to_assign_stmt_1351/type_cast_1337_Update/$entry
      -- CP-element group 420: 	 branch_block_stmt_33/assign_stmt_1322_to_assign_stmt_1351/type_cast_1337_Sample/rr
      -- CP-element group 420: 	 branch_block_stmt_33/assign_stmt_1322_to_assign_stmt_1351/type_cast_1337_Sample/$entry
      -- CP-element group 420: 	 branch_block_stmt_33/assign_stmt_1322_to_assign_stmt_1351/type_cast_1337_update_start_
      -- CP-element group 420: 	 branch_block_stmt_33/assign_stmt_1322_to_assign_stmt_1351/type_cast_1337_sample_start_
      -- CP-element group 420: 	 branch_block_stmt_33/assign_stmt_1322_to_assign_stmt_1351/$entry
      -- CP-element group 420: 	 branch_block_stmt_33/if_stmt_1310_if_link/if_choice_transition
      -- CP-element group 420: 	 branch_block_stmt_33/if_stmt_1310_if_link/$exit
      -- CP-element group 420: 	 branch_block_stmt_33/forx_xend273_bbx_xnph
      -- CP-element group 420: 	 branch_block_stmt_33/forx_xend273_bbx_xnph_PhiReq/$entry
      -- CP-element group 420: 	 branch_block_stmt_33/forx_xend273_bbx_xnph_PhiReq/$exit
      -- CP-element group 420: 	 branch_block_stmt_33/merge_stmt_1316_PhiReqMerge
      -- CP-element group 420: 	 branch_block_stmt_33/merge_stmt_1316_PhiAck/$entry
      -- CP-element group 420: 	 branch_block_stmt_33/merge_stmt_1316_PhiAck/$exit
      -- CP-element group 420: 	 branch_block_stmt_33/merge_stmt_1316_PhiAck/dummy
      -- 
    if_choice_transition_3095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 420_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1310_branch_ack_1, ack => convTranspose_CP_39_elements(420)); -- 
    cr_3117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(420), ack => type_cast_1337_inst_req_1); -- 
    rr_3112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(420), ack => type_cast_1337_inst_req_0); -- 
    -- CP-element group 421:  transition  place  input  bypass 
    -- CP-element group 421: predecessors 
    -- CP-element group 421: 	419 
    -- CP-element group 421: successors 
    -- CP-element group 421: 	499 
    -- CP-element group 421:  members (5) 
      -- CP-element group 421: 	 branch_block_stmt_33/forx_xend273_forx_xend501
      -- CP-element group 421: 	 branch_block_stmt_33/if_stmt_1310_else_link/else_choice_transition
      -- CP-element group 421: 	 branch_block_stmt_33/if_stmt_1310_else_link/$exit
      -- CP-element group 421: 	 branch_block_stmt_33/forx_xend273_forx_xend501_PhiReq/$entry
      -- CP-element group 421: 	 branch_block_stmt_33/forx_xend273_forx_xend501_PhiReq/$exit
      -- 
    else_choice_transition_3099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 421_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1310_branch_ack_0, ack => convTranspose_CP_39_elements(421)); -- 
    -- CP-element group 422:  transition  input  bypass 
    -- CP-element group 422: predecessors 
    -- CP-element group 422: 	420 
    -- CP-element group 422: successors 
    -- CP-element group 422:  members (3) 
      -- CP-element group 422: 	 branch_block_stmt_33/assign_stmt_1322_to_assign_stmt_1351/type_cast_1337_Sample/ra
      -- CP-element group 422: 	 branch_block_stmt_33/assign_stmt_1322_to_assign_stmt_1351/type_cast_1337_Sample/$exit
      -- CP-element group 422: 	 branch_block_stmt_33/assign_stmt_1322_to_assign_stmt_1351/type_cast_1337_sample_completed_
      -- 
    ra_3113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 422_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1337_inst_ack_0, ack => convTranspose_CP_39_elements(422)); -- 
    -- CP-element group 423:  transition  place  input  bypass 
    -- CP-element group 423: predecessors 
    -- CP-element group 423: 	420 
    -- CP-element group 423: successors 
    -- CP-element group 423: 	493 
    -- CP-element group 423:  members (9) 
      -- CP-element group 423: 	 branch_block_stmt_33/assign_stmt_1322_to_assign_stmt_1351__exit__
      -- CP-element group 423: 	 branch_block_stmt_33/bbx_xnph_forx_xbody428
      -- CP-element group 423: 	 branch_block_stmt_33/assign_stmt_1322_to_assign_stmt_1351/type_cast_1337_Update/ca
      -- CP-element group 423: 	 branch_block_stmt_33/assign_stmt_1322_to_assign_stmt_1351/type_cast_1337_Update/$exit
      -- CP-element group 423: 	 branch_block_stmt_33/assign_stmt_1322_to_assign_stmt_1351/type_cast_1337_update_completed_
      -- CP-element group 423: 	 branch_block_stmt_33/assign_stmt_1322_to_assign_stmt_1351/$exit
      -- CP-element group 423: 	 branch_block_stmt_33/bbx_xnph_forx_xbody428_PhiReq/$entry
      -- CP-element group 423: 	 branch_block_stmt_33/bbx_xnph_forx_xbody428_PhiReq/phi_stmt_1354/$entry
      -- CP-element group 423: 	 branch_block_stmt_33/bbx_xnph_forx_xbody428_PhiReq/phi_stmt_1354/phi_stmt_1354_sources/$entry
      -- 
    ca_3118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 423_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1337_inst_ack_1, ack => convTranspose_CP_39_elements(423)); -- 
    -- CP-element group 424:  transition  input  bypass 
    -- CP-element group 424: predecessors 
    -- CP-element group 424: 	498 
    -- CP-element group 424: successors 
    -- CP-element group 424: 	469 
    -- CP-element group 424:  members (3) 
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/array_obj_ref_1366_final_index_sum_regn_sample_complete
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/array_obj_ref_1366_final_index_sum_regn_Sample/$exit
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/array_obj_ref_1366_final_index_sum_regn_Sample/ack
      -- 
    ack_3147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 424_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1366_index_offset_ack_0, ack => convTranspose_CP_39_elements(424)); -- 
    -- CP-element group 425:  transition  input  output  bypass 
    -- CP-element group 425: predecessors 
    -- CP-element group 425: 	498 
    -- CP-element group 425: successors 
    -- CP-element group 425: 	426 
    -- CP-element group 425:  members (11) 
      -- CP-element group 425: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/addr_of_1367_request/req
      -- CP-element group 425: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/array_obj_ref_1366_offset_calculated
      -- CP-element group 425: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/array_obj_ref_1366_final_index_sum_regn_Update/$exit
      -- CP-element group 425: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/array_obj_ref_1366_final_index_sum_regn_Update/ack
      -- CP-element group 425: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/array_obj_ref_1366_base_plus_offset/$entry
      -- CP-element group 425: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/array_obj_ref_1366_base_plus_offset/$exit
      -- CP-element group 425: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/array_obj_ref_1366_base_plus_offset/sum_rename_req
      -- CP-element group 425: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/array_obj_ref_1366_base_plus_offset/sum_rename_ack
      -- CP-element group 425: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/addr_of_1367_request/$entry
      -- CP-element group 425: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/array_obj_ref_1366_root_address_calculated
      -- CP-element group 425: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/addr_of_1367_sample_start_
      -- 
    ack_3152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 425_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1366_index_offset_ack_1, ack => convTranspose_CP_39_elements(425)); -- 
    req_3161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(425), ack => addr_of_1367_final_reg_req_0); -- 
    -- CP-element group 426:  transition  input  bypass 
    -- CP-element group 426: predecessors 
    -- CP-element group 426: 	425 
    -- CP-element group 426: successors 
    -- CP-element group 426:  members (3) 
      -- CP-element group 426: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/addr_of_1367_request/$exit
      -- CP-element group 426: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/addr_of_1367_request/ack
      -- CP-element group 426: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/addr_of_1367_sample_completed_
      -- 
    ack_3162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 426_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1367_final_reg_ack_0, ack => convTranspose_CP_39_elements(426)); -- 
    -- CP-element group 427:  join  fork  transition  input  output  bypass 
    -- CP-element group 427: predecessors 
    -- CP-element group 427: 	498 
    -- CP-element group 427: successors 
    -- CP-element group 427: 	428 
    -- CP-element group 427:  members (24) 
      -- CP-element group 427: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/addr_of_1367_complete/$exit
      -- CP-element group 427: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/addr_of_1367_complete/ack
      -- CP-element group 427: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/ptr_deref_1371_sample_start_
      -- CP-element group 427: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/addr_of_1367_update_completed_
      -- CP-element group 427: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/ptr_deref_1371_Sample/word_access_start/word_0/rr
      -- CP-element group 427: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/ptr_deref_1371_Sample/word_access_start/word_0/$entry
      -- CP-element group 427: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/ptr_deref_1371_Sample/word_access_start/$entry
      -- CP-element group 427: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/ptr_deref_1371_Sample/$entry
      -- CP-element group 427: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/ptr_deref_1371_word_addrgen/root_register_ack
      -- CP-element group 427: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/ptr_deref_1371_word_addrgen/root_register_req
      -- CP-element group 427: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/ptr_deref_1371_word_addrgen/$exit
      -- CP-element group 427: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/ptr_deref_1371_word_addrgen/$entry
      -- CP-element group 427: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/ptr_deref_1371_base_plus_offset/sum_rename_ack
      -- CP-element group 427: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/ptr_deref_1371_base_plus_offset/sum_rename_req
      -- CP-element group 427: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/ptr_deref_1371_base_plus_offset/$exit
      -- CP-element group 427: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/ptr_deref_1371_base_plus_offset/$entry
      -- CP-element group 427: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/ptr_deref_1371_base_addr_resize/base_resize_ack
      -- CP-element group 427: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/ptr_deref_1371_base_addr_resize/base_resize_req
      -- CP-element group 427: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/ptr_deref_1371_base_addr_resize/$exit
      -- CP-element group 427: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/ptr_deref_1371_base_addr_resize/$entry
      -- CP-element group 427: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/ptr_deref_1371_base_address_resized
      -- CP-element group 427: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/ptr_deref_1371_root_address_calculated
      -- CP-element group 427: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/ptr_deref_1371_word_address_calculated
      -- CP-element group 427: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/ptr_deref_1371_base_address_calculated
      -- 
    ack_3167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 427_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1367_final_reg_ack_1, ack => convTranspose_CP_39_elements(427)); -- 
    rr_3200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(427), ack => ptr_deref_1371_load_0_req_0); -- 
    -- CP-element group 428:  transition  input  bypass 
    -- CP-element group 428: predecessors 
    -- CP-element group 428: 	427 
    -- CP-element group 428: successors 
    -- CP-element group 428:  members (5) 
      -- CP-element group 428: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/ptr_deref_1371_sample_completed_
      -- CP-element group 428: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/ptr_deref_1371_Sample/word_access_start/word_0/ra
      -- CP-element group 428: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/ptr_deref_1371_Sample/word_access_start/word_0/$exit
      -- CP-element group 428: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/ptr_deref_1371_Sample/word_access_start/$exit
      -- CP-element group 428: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/ptr_deref_1371_Sample/$exit
      -- 
    ra_3201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 428_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1371_load_0_ack_0, ack => convTranspose_CP_39_elements(428)); -- 
    -- CP-element group 429:  fork  transition  input  output  bypass 
    -- CP-element group 429: predecessors 
    -- CP-element group 429: 	498 
    -- CP-element group 429: successors 
    -- CP-element group 429: 	430 
    -- CP-element group 429: 	432 
    -- CP-element group 429: 	434 
    -- CP-element group 429: 	436 
    -- CP-element group 429: 	438 
    -- CP-element group 429: 	440 
    -- CP-element group 429: 	442 
    -- CP-element group 429: 	444 
    -- CP-element group 429:  members (33) 
      -- CP-element group 429: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1425_Sample/$entry
      -- CP-element group 429: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1405_sample_start_
      -- CP-element group 429: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1425_Sample/rr
      -- CP-element group 429: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1435_Sample/$entry
      -- CP-element group 429: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1375_Sample/rr
      -- CP-element group 429: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1395_Sample/rr
      -- CP-element group 429: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1405_Sample/$entry
      -- CP-element group 429: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1435_sample_start_
      -- CP-element group 429: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1405_Sample/rr
      -- CP-element group 429: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1445_Sample/$entry
      -- CP-element group 429: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1445_Sample/rr
      -- CP-element group 429: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1385_sample_start_
      -- CP-element group 429: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1445_sample_start_
      -- CP-element group 429: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1375_Sample/$entry
      -- CP-element group 429: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1395_Sample/$entry
      -- CP-element group 429: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1375_sample_start_
      -- CP-element group 429: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1395_sample_start_
      -- CP-element group 429: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/ptr_deref_1371_Update/ptr_deref_1371_Merge/merge_ack
      -- CP-element group 429: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/ptr_deref_1371_Update/ptr_deref_1371_Merge/merge_req
      -- CP-element group 429: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/ptr_deref_1371_Update/ptr_deref_1371_Merge/$exit
      -- CP-element group 429: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/ptr_deref_1371_Update/ptr_deref_1371_Merge/$entry
      -- CP-element group 429: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/ptr_deref_1371_Update/word_access_complete/word_0/ca
      -- CP-element group 429: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1425_sample_start_
      -- CP-element group 429: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/ptr_deref_1371_Update/word_access_complete/word_0/$exit
      -- CP-element group 429: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1385_Sample/rr
      -- CP-element group 429: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/ptr_deref_1371_Update/word_access_complete/$exit
      -- CP-element group 429: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/ptr_deref_1371_Update/$exit
      -- CP-element group 429: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1415_Sample/rr
      -- CP-element group 429: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1415_Sample/$entry
      -- CP-element group 429: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1385_Sample/$entry
      -- CP-element group 429: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1435_Sample/rr
      -- CP-element group 429: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1415_sample_start_
      -- CP-element group 429: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/ptr_deref_1371_update_completed_
      -- 
    ca_3212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 429_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1371_load_0_ack_1, ack => convTranspose_CP_39_elements(429)); -- 
    rr_3225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(429), ack => type_cast_1375_inst_req_0); -- 
    rr_3239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(429), ack => type_cast_1385_inst_req_0); -- 
    rr_3253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(429), ack => type_cast_1395_inst_req_0); -- 
    rr_3267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(429), ack => type_cast_1405_inst_req_0); -- 
    rr_3281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(429), ack => type_cast_1415_inst_req_0); -- 
    rr_3295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(429), ack => type_cast_1425_inst_req_0); -- 
    rr_3309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(429), ack => type_cast_1435_inst_req_0); -- 
    rr_3323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(429), ack => type_cast_1445_inst_req_0); -- 
    -- CP-element group 430:  transition  input  bypass 
    -- CP-element group 430: predecessors 
    -- CP-element group 430: 	429 
    -- CP-element group 430: successors 
    -- CP-element group 430:  members (3) 
      -- CP-element group 430: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1375_Sample/$exit
      -- CP-element group 430: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1375_Sample/ra
      -- CP-element group 430: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1375_sample_completed_
      -- 
    ra_3226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 430_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1375_inst_ack_0, ack => convTranspose_CP_39_elements(430)); -- 
    -- CP-element group 431:  transition  input  bypass 
    -- CP-element group 431: predecessors 
    -- CP-element group 431: 	498 
    -- CP-element group 431: successors 
    -- CP-element group 431: 	466 
    -- CP-element group 431:  members (3) 
      -- CP-element group 431: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1375_Update/$exit
      -- CP-element group 431: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1375_Update/ca
      -- CP-element group 431: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1375_update_completed_
      -- 
    ca_3231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 431_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1375_inst_ack_1, ack => convTranspose_CP_39_elements(431)); -- 
    -- CP-element group 432:  transition  input  bypass 
    -- CP-element group 432: predecessors 
    -- CP-element group 432: 	429 
    -- CP-element group 432: successors 
    -- CP-element group 432:  members (3) 
      -- CP-element group 432: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1385_Sample/ra
      -- CP-element group 432: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1385_Sample/$exit
      -- CP-element group 432: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1385_sample_completed_
      -- 
    ra_3240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 432_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1385_inst_ack_0, ack => convTranspose_CP_39_elements(432)); -- 
    -- CP-element group 433:  transition  input  bypass 
    -- CP-element group 433: predecessors 
    -- CP-element group 433: 	498 
    -- CP-element group 433: successors 
    -- CP-element group 433: 	463 
    -- CP-element group 433:  members (3) 
      -- CP-element group 433: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1385_Update/ca
      -- CP-element group 433: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1385_Update/$exit
      -- CP-element group 433: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1385_update_completed_
      -- 
    ca_3245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 433_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1385_inst_ack_1, ack => convTranspose_CP_39_elements(433)); -- 
    -- CP-element group 434:  transition  input  bypass 
    -- CP-element group 434: predecessors 
    -- CP-element group 434: 	429 
    -- CP-element group 434: successors 
    -- CP-element group 434:  members (3) 
      -- CP-element group 434: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1395_Sample/$exit
      -- CP-element group 434: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1395_Sample/ra
      -- CP-element group 434: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1395_sample_completed_
      -- 
    ra_3254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 434_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1395_inst_ack_0, ack => convTranspose_CP_39_elements(434)); -- 
    -- CP-element group 435:  transition  input  bypass 
    -- CP-element group 435: predecessors 
    -- CP-element group 435: 	498 
    -- CP-element group 435: successors 
    -- CP-element group 435: 	460 
    -- CP-element group 435:  members (3) 
      -- CP-element group 435: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1395_Update/ca
      -- CP-element group 435: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1395_Update/$exit
      -- CP-element group 435: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1395_update_completed_
      -- 
    ca_3259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 435_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1395_inst_ack_1, ack => convTranspose_CP_39_elements(435)); -- 
    -- CP-element group 436:  transition  input  bypass 
    -- CP-element group 436: predecessors 
    -- CP-element group 436: 	429 
    -- CP-element group 436: successors 
    -- CP-element group 436:  members (3) 
      -- CP-element group 436: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1405_sample_completed_
      -- CP-element group 436: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1405_Sample/$exit
      -- CP-element group 436: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1405_Sample/ra
      -- 
    ra_3268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 436_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1405_inst_ack_0, ack => convTranspose_CP_39_elements(436)); -- 
    -- CP-element group 437:  transition  input  bypass 
    -- CP-element group 437: predecessors 
    -- CP-element group 437: 	498 
    -- CP-element group 437: successors 
    -- CP-element group 437: 	457 
    -- CP-element group 437:  members (3) 
      -- CP-element group 437: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1405_update_completed_
      -- CP-element group 437: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1405_Update/ca
      -- CP-element group 437: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1405_Update/$exit
      -- 
    ca_3273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 437_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1405_inst_ack_1, ack => convTranspose_CP_39_elements(437)); -- 
    -- CP-element group 438:  transition  input  bypass 
    -- CP-element group 438: predecessors 
    -- CP-element group 438: 	429 
    -- CP-element group 438: successors 
    -- CP-element group 438:  members (3) 
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1415_Sample/ra
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1415_Sample/$exit
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1415_sample_completed_
      -- 
    ra_3282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 438_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1415_inst_ack_0, ack => convTranspose_CP_39_elements(438)); -- 
    -- CP-element group 439:  transition  input  bypass 
    -- CP-element group 439: predecessors 
    -- CP-element group 439: 	498 
    -- CP-element group 439: successors 
    -- CP-element group 439: 	454 
    -- CP-element group 439:  members (3) 
      -- CP-element group 439: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1415_Update/ca
      -- CP-element group 439: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1415_Update/$exit
      -- CP-element group 439: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1415_update_completed_
      -- 
    ca_3287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 439_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1415_inst_ack_1, ack => convTranspose_CP_39_elements(439)); -- 
    -- CP-element group 440:  transition  input  bypass 
    -- CP-element group 440: predecessors 
    -- CP-element group 440: 	429 
    -- CP-element group 440: successors 
    -- CP-element group 440:  members (3) 
      -- CP-element group 440: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1425_Sample/ra
      -- CP-element group 440: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1425_Sample/$exit
      -- CP-element group 440: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1425_sample_completed_
      -- 
    ra_3296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 440_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1425_inst_ack_0, ack => convTranspose_CP_39_elements(440)); -- 
    -- CP-element group 441:  transition  input  bypass 
    -- CP-element group 441: predecessors 
    -- CP-element group 441: 	498 
    -- CP-element group 441: successors 
    -- CP-element group 441: 	451 
    -- CP-element group 441:  members (3) 
      -- CP-element group 441: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1425_Update/ca
      -- CP-element group 441: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1425_update_completed_
      -- CP-element group 441: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1425_Update/$exit
      -- 
    ca_3301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 441_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1425_inst_ack_1, ack => convTranspose_CP_39_elements(441)); -- 
    -- CP-element group 442:  transition  input  bypass 
    -- CP-element group 442: predecessors 
    -- CP-element group 442: 	429 
    -- CP-element group 442: successors 
    -- CP-element group 442:  members (3) 
      -- CP-element group 442: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1435_sample_completed_
      -- CP-element group 442: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1435_Sample/ra
      -- CP-element group 442: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1435_Sample/$exit
      -- 
    ra_3310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 442_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1435_inst_ack_0, ack => convTranspose_CP_39_elements(442)); -- 
    -- CP-element group 443:  transition  input  bypass 
    -- CP-element group 443: predecessors 
    -- CP-element group 443: 	498 
    -- CP-element group 443: successors 
    -- CP-element group 443: 	448 
    -- CP-element group 443:  members (3) 
      -- CP-element group 443: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1435_Update/ca
      -- CP-element group 443: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1435_Update/$exit
      -- CP-element group 443: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1435_update_completed_
      -- 
    ca_3315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 443_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1435_inst_ack_1, ack => convTranspose_CP_39_elements(443)); -- 
    -- CP-element group 444:  transition  input  bypass 
    -- CP-element group 444: predecessors 
    -- CP-element group 444: 	429 
    -- CP-element group 444: successors 
    -- CP-element group 444:  members (3) 
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1445_sample_completed_
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1445_Sample/$exit
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1445_Sample/ra
      -- 
    ra_3324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 444_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1445_inst_ack_0, ack => convTranspose_CP_39_elements(444)); -- 
    -- CP-element group 445:  transition  input  output  bypass 
    -- CP-element group 445: predecessors 
    -- CP-element group 445: 	498 
    -- CP-element group 445: successors 
    -- CP-element group 445: 	446 
    -- CP-element group 445:  members (6) 
      -- CP-element group 445: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1445_update_completed_
      -- CP-element group 445: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1447_Sample/req
      -- CP-element group 445: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1447_Sample/$entry
      -- CP-element group 445: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1447_sample_start_
      -- CP-element group 445: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1445_Update/ca
      -- CP-element group 445: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1445_Update/$exit
      -- 
    ca_3329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 445_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1445_inst_ack_1, ack => convTranspose_CP_39_elements(445)); -- 
    req_3337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(445), ack => WPIPE_ConvTranspose_output_pipe_1447_inst_req_0); -- 
    -- CP-element group 446:  transition  input  output  bypass 
    -- CP-element group 446: predecessors 
    -- CP-element group 446: 	445 
    -- CP-element group 446: successors 
    -- CP-element group 446: 	447 
    -- CP-element group 446:  members (6) 
      -- CP-element group 446: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1447_Update/req
      -- CP-element group 446: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1447_Update/$entry
      -- CP-element group 446: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1447_Sample/ack
      -- CP-element group 446: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1447_Sample/$exit
      -- CP-element group 446: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1447_update_start_
      -- CP-element group 446: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1447_sample_completed_
      -- 
    ack_3338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 446_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1447_inst_ack_0, ack => convTranspose_CP_39_elements(446)); -- 
    req_3342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(446), ack => WPIPE_ConvTranspose_output_pipe_1447_inst_req_1); -- 
    -- CP-element group 447:  transition  input  bypass 
    -- CP-element group 447: predecessors 
    -- CP-element group 447: 	446 
    -- CP-element group 447: successors 
    -- CP-element group 447: 	448 
    -- CP-element group 447:  members (3) 
      -- CP-element group 447: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1447_Update/ack
      -- CP-element group 447: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1447_Update/$exit
      -- CP-element group 447: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1447_update_completed_
      -- 
    ack_3343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 447_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1447_inst_ack_1, ack => convTranspose_CP_39_elements(447)); -- 
    -- CP-element group 448:  join  transition  output  bypass 
    -- CP-element group 448: predecessors 
    -- CP-element group 448: 	443 
    -- CP-element group 448: 	447 
    -- CP-element group 448: successors 
    -- CP-element group 448: 	449 
    -- CP-element group 448:  members (3) 
      -- CP-element group 448: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1450_Sample/req
      -- CP-element group 448: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1450_Sample/$entry
      -- CP-element group 448: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1450_sample_start_
      -- 
    req_3351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(448), ack => WPIPE_ConvTranspose_output_pipe_1450_inst_req_0); -- 
    convTranspose_cp_element_group_448: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_448"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(443) & convTranspose_CP_39_elements(447);
      gj_convTranspose_cp_element_group_448 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(448), clk => clk, reset => reset); --
    end block;
    -- CP-element group 449:  transition  input  output  bypass 
    -- CP-element group 449: predecessors 
    -- CP-element group 449: 	448 
    -- CP-element group 449: successors 
    -- CP-element group 449: 	450 
    -- CP-element group 449:  members (6) 
      -- CP-element group 449: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1450_Update/req
      -- CP-element group 449: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1450_Update/$entry
      -- CP-element group 449: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1450_Sample/ack
      -- CP-element group 449: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1450_Sample/$exit
      -- CP-element group 449: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1450_update_start_
      -- CP-element group 449: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1450_sample_completed_
      -- 
    ack_3352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 449_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1450_inst_ack_0, ack => convTranspose_CP_39_elements(449)); -- 
    req_3356_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3356_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(449), ack => WPIPE_ConvTranspose_output_pipe_1450_inst_req_1); -- 
    -- CP-element group 450:  transition  input  bypass 
    -- CP-element group 450: predecessors 
    -- CP-element group 450: 	449 
    -- CP-element group 450: successors 
    -- CP-element group 450: 	451 
    -- CP-element group 450:  members (3) 
      -- CP-element group 450: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1450_Update/ack
      -- CP-element group 450: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1450_Update/$exit
      -- CP-element group 450: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1450_update_completed_
      -- 
    ack_3357_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 450_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1450_inst_ack_1, ack => convTranspose_CP_39_elements(450)); -- 
    -- CP-element group 451:  join  transition  output  bypass 
    -- CP-element group 451: predecessors 
    -- CP-element group 451: 	441 
    -- CP-element group 451: 	450 
    -- CP-element group 451: successors 
    -- CP-element group 451: 	452 
    -- CP-element group 451:  members (3) 
      -- CP-element group 451: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1453_Sample/$entry
      -- CP-element group 451: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1453_sample_start_
      -- CP-element group 451: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1453_Sample/req
      -- 
    req_3365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(451), ack => WPIPE_ConvTranspose_output_pipe_1453_inst_req_0); -- 
    convTranspose_cp_element_group_451: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_451"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(441) & convTranspose_CP_39_elements(450);
      gj_convTranspose_cp_element_group_451 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(451), clk => clk, reset => reset); --
    end block;
    -- CP-element group 452:  transition  input  output  bypass 
    -- CP-element group 452: predecessors 
    -- CP-element group 452: 	451 
    -- CP-element group 452: successors 
    -- CP-element group 452: 	453 
    -- CP-element group 452:  members (6) 
      -- CP-element group 452: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1453_Sample/$exit
      -- CP-element group 452: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1453_update_start_
      -- CP-element group 452: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1453_sample_completed_
      -- CP-element group 452: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1453_Update/req
      -- CP-element group 452: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1453_Update/$entry
      -- CP-element group 452: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1453_Sample/ack
      -- 
    ack_3366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 452_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1453_inst_ack_0, ack => convTranspose_CP_39_elements(452)); -- 
    req_3370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(452), ack => WPIPE_ConvTranspose_output_pipe_1453_inst_req_1); -- 
    -- CP-element group 453:  transition  input  bypass 
    -- CP-element group 453: predecessors 
    -- CP-element group 453: 	452 
    -- CP-element group 453: successors 
    -- CP-element group 453: 	454 
    -- CP-element group 453:  members (3) 
      -- CP-element group 453: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1453_update_completed_
      -- CP-element group 453: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1453_Update/ack
      -- CP-element group 453: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1453_Update/$exit
      -- 
    ack_3371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 453_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1453_inst_ack_1, ack => convTranspose_CP_39_elements(453)); -- 
    -- CP-element group 454:  join  transition  output  bypass 
    -- CP-element group 454: predecessors 
    -- CP-element group 454: 	439 
    -- CP-element group 454: 	453 
    -- CP-element group 454: successors 
    -- CP-element group 454: 	455 
    -- CP-element group 454:  members (3) 
      -- CP-element group 454: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1456_sample_start_
      -- CP-element group 454: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1456_Sample/$entry
      -- CP-element group 454: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1456_Sample/req
      -- 
    req_3379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(454), ack => WPIPE_ConvTranspose_output_pipe_1456_inst_req_0); -- 
    convTranspose_cp_element_group_454: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_454"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(439) & convTranspose_CP_39_elements(453);
      gj_convTranspose_cp_element_group_454 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(454), clk => clk, reset => reset); --
    end block;
    -- CP-element group 455:  transition  input  output  bypass 
    -- CP-element group 455: predecessors 
    -- CP-element group 455: 	454 
    -- CP-element group 455: successors 
    -- CP-element group 455: 	456 
    -- CP-element group 455:  members (6) 
      -- CP-element group 455: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1456_sample_completed_
      -- CP-element group 455: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1456_update_start_
      -- CP-element group 455: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1456_Sample/$exit
      -- CP-element group 455: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1456_Sample/ack
      -- CP-element group 455: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1456_Update/$entry
      -- CP-element group 455: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1456_Update/req
      -- 
    ack_3380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 455_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1456_inst_ack_0, ack => convTranspose_CP_39_elements(455)); -- 
    req_3384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(455), ack => WPIPE_ConvTranspose_output_pipe_1456_inst_req_1); -- 
    -- CP-element group 456:  transition  input  bypass 
    -- CP-element group 456: predecessors 
    -- CP-element group 456: 	455 
    -- CP-element group 456: successors 
    -- CP-element group 456: 	457 
    -- CP-element group 456:  members (3) 
      -- CP-element group 456: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1456_update_completed_
      -- CP-element group 456: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1456_Update/$exit
      -- CP-element group 456: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1456_Update/ack
      -- 
    ack_3385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 456_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1456_inst_ack_1, ack => convTranspose_CP_39_elements(456)); -- 
    -- CP-element group 457:  join  transition  output  bypass 
    -- CP-element group 457: predecessors 
    -- CP-element group 457: 	437 
    -- CP-element group 457: 	456 
    -- CP-element group 457: successors 
    -- CP-element group 457: 	458 
    -- CP-element group 457:  members (3) 
      -- CP-element group 457: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1459_sample_start_
      -- CP-element group 457: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1459_Sample/$entry
      -- CP-element group 457: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1459_Sample/req
      -- 
    req_3393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(457), ack => WPIPE_ConvTranspose_output_pipe_1459_inst_req_0); -- 
    convTranspose_cp_element_group_457: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_457"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(437) & convTranspose_CP_39_elements(456);
      gj_convTranspose_cp_element_group_457 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(457), clk => clk, reset => reset); --
    end block;
    -- CP-element group 458:  transition  input  output  bypass 
    -- CP-element group 458: predecessors 
    -- CP-element group 458: 	457 
    -- CP-element group 458: successors 
    -- CP-element group 458: 	459 
    -- CP-element group 458:  members (6) 
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1459_sample_completed_
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1459_update_start_
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1459_Sample/$exit
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1459_Sample/ack
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1459_Update/$entry
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1459_Update/req
      -- 
    ack_3394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 458_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1459_inst_ack_0, ack => convTranspose_CP_39_elements(458)); -- 
    req_3398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(458), ack => WPIPE_ConvTranspose_output_pipe_1459_inst_req_1); -- 
    -- CP-element group 459:  transition  input  bypass 
    -- CP-element group 459: predecessors 
    -- CP-element group 459: 	458 
    -- CP-element group 459: successors 
    -- CP-element group 459: 	460 
    -- CP-element group 459:  members (3) 
      -- CP-element group 459: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1459_update_completed_
      -- CP-element group 459: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1459_Update/$exit
      -- CP-element group 459: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1459_Update/ack
      -- 
    ack_3399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 459_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1459_inst_ack_1, ack => convTranspose_CP_39_elements(459)); -- 
    -- CP-element group 460:  join  transition  output  bypass 
    -- CP-element group 460: predecessors 
    -- CP-element group 460: 	435 
    -- CP-element group 460: 	459 
    -- CP-element group 460: successors 
    -- CP-element group 460: 	461 
    -- CP-element group 460:  members (3) 
      -- CP-element group 460: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1462_sample_start_
      -- CP-element group 460: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1462_Sample/$entry
      -- CP-element group 460: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1462_Sample/req
      -- 
    req_3407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(460), ack => WPIPE_ConvTranspose_output_pipe_1462_inst_req_0); -- 
    convTranspose_cp_element_group_460: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_460"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(435) & convTranspose_CP_39_elements(459);
      gj_convTranspose_cp_element_group_460 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(460), clk => clk, reset => reset); --
    end block;
    -- CP-element group 461:  transition  input  output  bypass 
    -- CP-element group 461: predecessors 
    -- CP-element group 461: 	460 
    -- CP-element group 461: successors 
    -- CP-element group 461: 	462 
    -- CP-element group 461:  members (6) 
      -- CP-element group 461: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1462_sample_completed_
      -- CP-element group 461: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1462_update_start_
      -- CP-element group 461: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1462_Sample/$exit
      -- CP-element group 461: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1462_Sample/ack
      -- CP-element group 461: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1462_Update/$entry
      -- CP-element group 461: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1462_Update/req
      -- 
    ack_3408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 461_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1462_inst_ack_0, ack => convTranspose_CP_39_elements(461)); -- 
    req_3412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(461), ack => WPIPE_ConvTranspose_output_pipe_1462_inst_req_1); -- 
    -- CP-element group 462:  transition  input  bypass 
    -- CP-element group 462: predecessors 
    -- CP-element group 462: 	461 
    -- CP-element group 462: successors 
    -- CP-element group 462: 	463 
    -- CP-element group 462:  members (3) 
      -- CP-element group 462: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1462_update_completed_
      -- CP-element group 462: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1462_Update/$exit
      -- CP-element group 462: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1462_Update/ack
      -- 
    ack_3413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 462_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1462_inst_ack_1, ack => convTranspose_CP_39_elements(462)); -- 
    -- CP-element group 463:  join  transition  output  bypass 
    -- CP-element group 463: predecessors 
    -- CP-element group 463: 	433 
    -- CP-element group 463: 	462 
    -- CP-element group 463: successors 
    -- CP-element group 463: 	464 
    -- CP-element group 463:  members (3) 
      -- CP-element group 463: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1465_sample_start_
      -- CP-element group 463: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1465_Sample/$entry
      -- CP-element group 463: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1465_Sample/req
      -- 
    req_3421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(463), ack => WPIPE_ConvTranspose_output_pipe_1465_inst_req_0); -- 
    convTranspose_cp_element_group_463: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_463"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(433) & convTranspose_CP_39_elements(462);
      gj_convTranspose_cp_element_group_463 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(463), clk => clk, reset => reset); --
    end block;
    -- CP-element group 464:  transition  input  output  bypass 
    -- CP-element group 464: predecessors 
    -- CP-element group 464: 	463 
    -- CP-element group 464: successors 
    -- CP-element group 464: 	465 
    -- CP-element group 464:  members (6) 
      -- CP-element group 464: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1465_sample_completed_
      -- CP-element group 464: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1465_update_start_
      -- CP-element group 464: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1465_Sample/$exit
      -- CP-element group 464: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1465_Sample/ack
      -- CP-element group 464: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1465_Update/$entry
      -- CP-element group 464: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1465_Update/req
      -- 
    ack_3422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 464_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1465_inst_ack_0, ack => convTranspose_CP_39_elements(464)); -- 
    req_3426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(464), ack => WPIPE_ConvTranspose_output_pipe_1465_inst_req_1); -- 
    -- CP-element group 465:  transition  input  bypass 
    -- CP-element group 465: predecessors 
    -- CP-element group 465: 	464 
    -- CP-element group 465: successors 
    -- CP-element group 465: 	466 
    -- CP-element group 465:  members (3) 
      -- CP-element group 465: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1465_update_completed_
      -- CP-element group 465: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1465_Update/$exit
      -- CP-element group 465: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1465_Update/ack
      -- 
    ack_3427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 465_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1465_inst_ack_1, ack => convTranspose_CP_39_elements(465)); -- 
    -- CP-element group 466:  join  transition  output  bypass 
    -- CP-element group 466: predecessors 
    -- CP-element group 466: 	431 
    -- CP-element group 466: 	465 
    -- CP-element group 466: successors 
    -- CP-element group 466: 	467 
    -- CP-element group 466:  members (3) 
      -- CP-element group 466: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1468_sample_start_
      -- CP-element group 466: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1468_Sample/$entry
      -- CP-element group 466: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1468_Sample/req
      -- 
    req_3435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(466), ack => WPIPE_ConvTranspose_output_pipe_1468_inst_req_0); -- 
    convTranspose_cp_element_group_466: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_466"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(431) & convTranspose_CP_39_elements(465);
      gj_convTranspose_cp_element_group_466 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(466), clk => clk, reset => reset); --
    end block;
    -- CP-element group 467:  transition  input  output  bypass 
    -- CP-element group 467: predecessors 
    -- CP-element group 467: 	466 
    -- CP-element group 467: successors 
    -- CP-element group 467: 	468 
    -- CP-element group 467:  members (6) 
      -- CP-element group 467: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1468_sample_completed_
      -- CP-element group 467: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1468_update_start_
      -- CP-element group 467: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1468_Sample/$exit
      -- CP-element group 467: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1468_Sample/ack
      -- CP-element group 467: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1468_Update/$entry
      -- CP-element group 467: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1468_Update/req
      -- 
    ack_3436_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 467_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1468_inst_ack_0, ack => convTranspose_CP_39_elements(467)); -- 
    req_3440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(467), ack => WPIPE_ConvTranspose_output_pipe_1468_inst_req_1); -- 
    -- CP-element group 468:  transition  input  bypass 
    -- CP-element group 468: predecessors 
    -- CP-element group 468: 	467 
    -- CP-element group 468: successors 
    -- CP-element group 468: 	469 
    -- CP-element group 468:  members (3) 
      -- CP-element group 468: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1468_update_completed_
      -- CP-element group 468: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1468_Update/$exit
      -- CP-element group 468: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/WPIPE_ConvTranspose_output_pipe_1468_Update/ack
      -- 
    ack_3441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 468_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1468_inst_ack_1, ack => convTranspose_CP_39_elements(468)); -- 
    -- CP-element group 469:  branch  join  transition  place  output  bypass 
    -- CP-element group 469: predecessors 
    -- CP-element group 469: 	424 
    -- CP-element group 469: 	468 
    -- CP-element group 469: successors 
    -- CP-element group 469: 	470 
    -- CP-element group 469: 	471 
    -- CP-element group 469:  members (10) 
      -- CP-element group 469: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481__exit__
      -- CP-element group 469: 	 branch_block_stmt_33/if_stmt_1482__entry__
      -- CP-element group 469: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/$exit
      -- CP-element group 469: 	 branch_block_stmt_33/if_stmt_1482_dead_link/$entry
      -- CP-element group 469: 	 branch_block_stmt_33/if_stmt_1482_eval_test/$entry
      -- CP-element group 469: 	 branch_block_stmt_33/if_stmt_1482_eval_test/$exit
      -- CP-element group 469: 	 branch_block_stmt_33/if_stmt_1482_eval_test/branch_req
      -- CP-element group 469: 	 branch_block_stmt_33/R_exitcond1_1483_place
      -- CP-element group 469: 	 branch_block_stmt_33/if_stmt_1482_if_link/$entry
      -- CP-element group 469: 	 branch_block_stmt_33/if_stmt_1482_else_link/$entry
      -- 
    branch_req_3449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(469), ack => if_stmt_1482_branch_req_0); -- 
    convTranspose_cp_element_group_469: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_469"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(424) & convTranspose_CP_39_elements(468);
      gj_convTranspose_cp_element_group_469 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(469), clk => clk, reset => reset); --
    end block;
    -- CP-element group 470:  merge  transition  place  input  bypass 
    -- CP-element group 470: predecessors 
    -- CP-element group 470: 	469 
    -- CP-element group 470: successors 
    -- CP-element group 470: 	499 
    -- CP-element group 470:  members (13) 
      -- CP-element group 470: 	 branch_block_stmt_33/merge_stmt_1488__exit__
      -- CP-element group 470: 	 branch_block_stmt_33/forx_xend501x_xloopexit_forx_xend501
      -- CP-element group 470: 	 branch_block_stmt_33/if_stmt_1482_if_link/$exit
      -- CP-element group 470: 	 branch_block_stmt_33/if_stmt_1482_if_link/if_choice_transition
      -- CP-element group 470: 	 branch_block_stmt_33/forx_xbody428_forx_xend501x_xloopexit
      -- CP-element group 470: 	 branch_block_stmt_33/forx_xbody428_forx_xend501x_xloopexit_PhiReq/$entry
      -- CP-element group 470: 	 branch_block_stmt_33/forx_xbody428_forx_xend501x_xloopexit_PhiReq/$exit
      -- CP-element group 470: 	 branch_block_stmt_33/merge_stmt_1488_PhiReqMerge
      -- CP-element group 470: 	 branch_block_stmt_33/merge_stmt_1488_PhiAck/$entry
      -- CP-element group 470: 	 branch_block_stmt_33/merge_stmt_1488_PhiAck/$exit
      -- CP-element group 470: 	 branch_block_stmt_33/merge_stmt_1488_PhiAck/dummy
      -- CP-element group 470: 	 branch_block_stmt_33/forx_xend501x_xloopexit_forx_xend501_PhiReq/$entry
      -- CP-element group 470: 	 branch_block_stmt_33/forx_xend501x_xloopexit_forx_xend501_PhiReq/$exit
      -- 
    if_choice_transition_3454_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 470_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1482_branch_ack_1, ack => convTranspose_CP_39_elements(470)); -- 
    -- CP-element group 471:  fork  transition  place  input  output  bypass 
    -- CP-element group 471: predecessors 
    -- CP-element group 471: 	469 
    -- CP-element group 471: successors 
    -- CP-element group 471: 	494 
    -- CP-element group 471: 	495 
    -- CP-element group 471:  members (12) 
      -- CP-element group 471: 	 branch_block_stmt_33/if_stmt_1482_else_link/$exit
      -- CP-element group 471: 	 branch_block_stmt_33/if_stmt_1482_else_link/else_choice_transition
      -- CP-element group 471: 	 branch_block_stmt_33/forx_xbody428_forx_xbody428
      -- CP-element group 471: 	 branch_block_stmt_33/forx_xbody428_forx_xbody428_PhiReq/$entry
      -- CP-element group 471: 	 branch_block_stmt_33/forx_xbody428_forx_xbody428_PhiReq/phi_stmt_1354/$entry
      -- CP-element group 471: 	 branch_block_stmt_33/forx_xbody428_forx_xbody428_PhiReq/phi_stmt_1354/phi_stmt_1354_sources/$entry
      -- CP-element group 471: 	 branch_block_stmt_33/forx_xbody428_forx_xbody428_PhiReq/phi_stmt_1354/phi_stmt_1354_sources/type_cast_1360/$entry
      -- CP-element group 471: 	 branch_block_stmt_33/forx_xbody428_forx_xbody428_PhiReq/phi_stmt_1354/phi_stmt_1354_sources/type_cast_1360/SplitProtocol/$entry
      -- CP-element group 471: 	 branch_block_stmt_33/forx_xbody428_forx_xbody428_PhiReq/phi_stmt_1354/phi_stmt_1354_sources/type_cast_1360/SplitProtocol/Sample/$entry
      -- CP-element group 471: 	 branch_block_stmt_33/forx_xbody428_forx_xbody428_PhiReq/phi_stmt_1354/phi_stmt_1354_sources/type_cast_1360/SplitProtocol/Sample/rr
      -- CP-element group 471: 	 branch_block_stmt_33/forx_xbody428_forx_xbody428_PhiReq/phi_stmt_1354/phi_stmt_1354_sources/type_cast_1360/SplitProtocol/Update/$entry
      -- CP-element group 471: 	 branch_block_stmt_33/forx_xbody428_forx_xbody428_PhiReq/phi_stmt_1354/phi_stmt_1354_sources/type_cast_1360/SplitProtocol/Update/cr
      -- 
    else_choice_transition_3458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 471_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1482_branch_ack_0, ack => convTranspose_CP_39_elements(471)); -- 
    rr_3733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(471), ack => type_cast_1360_inst_req_0); -- 
    cr_3738_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3738_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(471), ack => type_cast_1360_inst_req_1); -- 
    -- CP-element group 472:  merge  branch  transition  place  output  bypass 
    -- CP-element group 472: predecessors 
    -- CP-element group 472: 	165 
    -- CP-element group 472: 	120 
    -- CP-element group 472: successors 
    -- CP-element group 472: 	121 
    -- CP-element group 472: 	122 
    -- CP-element group 472:  members (17) 
      -- CP-element group 472: 	 branch_block_stmt_33/merge_stmt_425__exit__
      -- CP-element group 472: 	 branch_block_stmt_33/assign_stmt_431__entry__
      -- CP-element group 472: 	 branch_block_stmt_33/assign_stmt_431__exit__
      -- CP-element group 472: 	 branch_block_stmt_33/if_stmt_432__entry__
      -- CP-element group 472: 	 branch_block_stmt_33/assign_stmt_431/$entry
      -- CP-element group 472: 	 branch_block_stmt_33/assign_stmt_431/$exit
      -- CP-element group 472: 	 branch_block_stmt_33/if_stmt_432_dead_link/$entry
      -- CP-element group 472: 	 branch_block_stmt_33/if_stmt_432_eval_test/$entry
      -- CP-element group 472: 	 branch_block_stmt_33/if_stmt_432_eval_test/$exit
      -- CP-element group 472: 	 branch_block_stmt_33/if_stmt_432_eval_test/branch_req
      -- CP-element group 472: 	 branch_block_stmt_33/R_cmp194510_433_place
      -- CP-element group 472: 	 branch_block_stmt_33/if_stmt_432_if_link/$entry
      -- CP-element group 472: 	 branch_block_stmt_33/if_stmt_432_else_link/$entry
      -- CP-element group 472: 	 branch_block_stmt_33/merge_stmt_425_PhiReqMerge
      -- CP-element group 472: 	 branch_block_stmt_33/merge_stmt_425_PhiAck/$entry
      -- CP-element group 472: 	 branch_block_stmt_33/merge_stmt_425_PhiAck/$exit
      -- CP-element group 472: 	 branch_block_stmt_33/merge_stmt_425_PhiAck/dummy
      -- 
    branch_req_927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(472), ack => if_stmt_432_branch_req_0); -- 
    convTranspose_CP_39_elements(472) <= OrReduce(convTranspose_CP_39_elements(165) & convTranspose_CP_39_elements(120));
    -- CP-element group 473:  transition  output  delay-element  bypass 
    -- CP-element group 473: predecessors 
    -- CP-element group 473: 	124 
    -- CP-element group 473: successors 
    -- CP-element group 473: 	477 
    -- CP-element group 473:  members (5) 
      -- CP-element group 473: 	 branch_block_stmt_33/bbx_xnph516_forx_xbody_PhiReq/$exit
      -- CP-element group 473: 	 branch_block_stmt_33/bbx_xnph516_forx_xbody_PhiReq/phi_stmt_470/$exit
      -- CP-element group 473: 	 branch_block_stmt_33/bbx_xnph516_forx_xbody_PhiReq/phi_stmt_470/phi_stmt_470_sources/$exit
      -- CP-element group 473: 	 branch_block_stmt_33/bbx_xnph516_forx_xbody_PhiReq/phi_stmt_470/phi_stmt_470_sources/type_cast_474_konst_delay_trans
      -- CP-element group 473: 	 branch_block_stmt_33/bbx_xnph516_forx_xbody_PhiReq/phi_stmt_470/phi_stmt_470_req
      -- 
    phi_stmt_470_req_3506_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_470_req_3506_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(473), ack => phi_stmt_470_req_0); -- 
    -- Element group convTranspose_CP_39_elements(473) is a control-delay.
    cp_element_473_delay: control_delay_element  generic map(name => " 473_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(124), ack => convTranspose_CP_39_elements(473), clk => clk, reset =>reset);
    -- CP-element group 474:  transition  input  bypass 
    -- CP-element group 474: predecessors 
    -- CP-element group 474: 	166 
    -- CP-element group 474: successors 
    -- CP-element group 474: 	476 
    -- CP-element group 474:  members (2) 
      -- CP-element group 474: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_470/phi_stmt_470_sources/type_cast_476/SplitProtocol/Sample/$exit
      -- CP-element group 474: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_470/phi_stmt_470_sources/type_cast_476/SplitProtocol/Sample/ra
      -- 
    ra_3526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 474_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_476_inst_ack_0, ack => convTranspose_CP_39_elements(474)); -- 
    -- CP-element group 475:  transition  input  bypass 
    -- CP-element group 475: predecessors 
    -- CP-element group 475: 	166 
    -- CP-element group 475: successors 
    -- CP-element group 475: 	476 
    -- CP-element group 475:  members (2) 
      -- CP-element group 475: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_470/phi_stmt_470_sources/type_cast_476/SplitProtocol/Update/$exit
      -- CP-element group 475: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_470/phi_stmt_470_sources/type_cast_476/SplitProtocol/Update/ca
      -- 
    ca_3531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 475_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_476_inst_ack_1, ack => convTranspose_CP_39_elements(475)); -- 
    -- CP-element group 476:  join  transition  output  bypass 
    -- CP-element group 476: predecessors 
    -- CP-element group 476: 	474 
    -- CP-element group 476: 	475 
    -- CP-element group 476: successors 
    -- CP-element group 476: 	477 
    -- CP-element group 476:  members (6) 
      -- CP-element group 476: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 476: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_470/$exit
      -- CP-element group 476: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_470/phi_stmt_470_sources/$exit
      -- CP-element group 476: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_470/phi_stmt_470_sources/type_cast_476/$exit
      -- CP-element group 476: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_470/phi_stmt_470_sources/type_cast_476/SplitProtocol/$exit
      -- CP-element group 476: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_470/phi_stmt_470_req
      -- 
    phi_stmt_470_req_3532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_470_req_3532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(476), ack => phi_stmt_470_req_1); -- 
    convTranspose_cp_element_group_476: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_476"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(474) & convTranspose_CP_39_elements(475);
      gj_convTranspose_cp_element_group_476 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(476), clk => clk, reset => reset); --
    end block;
    -- CP-element group 477:  merge  transition  place  bypass 
    -- CP-element group 477: predecessors 
    -- CP-element group 477: 	473 
    -- CP-element group 477: 	476 
    -- CP-element group 477: successors 
    -- CP-element group 477: 	478 
    -- CP-element group 477:  members (2) 
      -- CP-element group 477: 	 branch_block_stmt_33/merge_stmt_469_PhiReqMerge
      -- CP-element group 477: 	 branch_block_stmt_33/merge_stmt_469_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(477) <= OrReduce(convTranspose_CP_39_elements(473) & convTranspose_CP_39_elements(476));
    -- CP-element group 478:  fork  transition  place  input  output  bypass 
    -- CP-element group 478: predecessors 
    -- CP-element group 478: 	477 
    -- CP-element group 478: successors 
    -- CP-element group 478: 	156 
    -- CP-element group 478: 	160 
    -- CP-element group 478: 	163 
    -- CP-element group 478: 	125 
    -- CP-element group 478: 	126 
    -- CP-element group 478: 	128 
    -- CP-element group 478: 	129 
    -- CP-element group 478: 	132 
    -- CP-element group 478: 	136 
    -- CP-element group 478: 	140 
    -- CP-element group 478: 	144 
    -- CP-element group 478: 	148 
    -- CP-element group 478: 	152 
    -- CP-element group 478:  members (56) 
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_611_update_start_
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_575_Update/cr
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_575_Update/$entry
      -- CP-element group 478: 	 branch_block_stmt_33/merge_stmt_469__exit__
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632__entry__
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_539_update_start_
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_575_update_start_
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_557_Update/cr
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_557_Update/$entry
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_521_Update/cr
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_557_update_start_
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_update_start_
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_Update/word_access_complete/word_0/cr
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_521_Update/$entry
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_Update/word_access_complete/word_0/$entry
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_593_Update/cr
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_Update/word_access_complete/$entry
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_593_Update/$entry
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_Update/$entry
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_611_Update/cr
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_611_Update/$entry
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_539_Update/cr
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_593_update_start_
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_539_Update/$entry
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/$entry
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/addr_of_483_update_start_
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_index_resized_1
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_index_scaled_1
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_index_computed_1
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_index_resize_1/$entry
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_index_resize_1/$exit
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_index_resize_1/index_resize_req
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_index_resize_1/index_resize_ack
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_index_scale_1/$entry
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_index_scale_1/$exit
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_index_scale_1/scale_rename_req
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_index_scale_1/scale_rename_ack
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_final_index_sum_regn_update_start
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_final_index_sum_regn_Sample/$entry
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_final_index_sum_regn_Sample/req
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_final_index_sum_regn_Update/$entry
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_final_index_sum_regn_Update/req
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/addr_of_483_complete/$entry
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/addr_of_483_complete/req
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_486_sample_start_
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_486_Sample/$entry
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_486_Sample/rr
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_490_update_start_
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_490_Update/$entry
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_490_Update/cr
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_503_update_start_
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_503_Update/$entry
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_503_Update/cr
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_521_update_start_
      -- CP-element group 478: 	 branch_block_stmt_33/merge_stmt_469_PhiAck/$exit
      -- CP-element group 478: 	 branch_block_stmt_33/merge_stmt_469_PhiAck/phi_stmt_470_ack
      -- 
    phi_stmt_470_ack_3537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 478_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_470_ack_0, ack => convTranspose_CP_39_elements(478)); -- 
    cr_1171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(478), ack => type_cast_575_inst_req_1); -- 
    cr_1143_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1143_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(478), ack => type_cast_557_inst_req_1); -- 
    cr_1087_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1087_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(478), ack => type_cast_521_inst_req_1); -- 
    cr_1277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(478), ack => ptr_deref_619_store_0_req_1); -- 
    cr_1199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(478), ack => type_cast_593_inst_req_1); -- 
    cr_1227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(478), ack => type_cast_611_inst_req_1); -- 
    cr_1115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(478), ack => type_cast_539_inst_req_1); -- 
    req_983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(478), ack => array_obj_ref_482_index_offset_req_0); -- 
    req_988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(478), ack => array_obj_ref_482_index_offset_req_1); -- 
    req_1003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(478), ack => addr_of_483_final_reg_req_1); -- 
    rr_1012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(478), ack => RPIPE_ConvTranspose_input_pipe_486_inst_req_0); -- 
    cr_1031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(478), ack => type_cast_490_inst_req_1); -- 
    cr_1059_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1059_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(478), ack => type_cast_503_inst_req_1); -- 
    -- CP-element group 479:  transition  output  delay-element  bypass 
    -- CP-element group 479: predecessors 
    -- CP-element group 479: 	168 
    -- CP-element group 479: successors 
    -- CP-element group 479: 	483 
    -- CP-element group 479:  members (5) 
      -- CP-element group 479: 	 branch_block_stmt_33/bbx_xnph512_forx_xbody196_PhiReq/$exit
      -- CP-element group 479: 	 branch_block_stmt_33/bbx_xnph512_forx_xbody196_PhiReq/phi_stmt_677/$exit
      -- CP-element group 479: 	 branch_block_stmt_33/bbx_xnph512_forx_xbody196_PhiReq/phi_stmt_677/phi_stmt_677_sources/$exit
      -- CP-element group 479: 	 branch_block_stmt_33/bbx_xnph512_forx_xbody196_PhiReq/phi_stmt_677/phi_stmt_677_sources/type_cast_681_konst_delay_trans
      -- CP-element group 479: 	 branch_block_stmt_33/bbx_xnph512_forx_xbody196_PhiReq/phi_stmt_677/phi_stmt_677_req
      -- 
    phi_stmt_677_req_3560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_677_req_3560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(479), ack => phi_stmt_677_req_0); -- 
    -- Element group convTranspose_CP_39_elements(479) is a control-delay.
    cp_element_479_delay: control_delay_element  generic map(name => " 479_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(168), ack => convTranspose_CP_39_elements(479), clk => clk, reset =>reset);
    -- CP-element group 480:  transition  input  bypass 
    -- CP-element group 480: predecessors 
    -- CP-element group 480: 	210 
    -- CP-element group 480: successors 
    -- CP-element group 480: 	482 
    -- CP-element group 480:  members (2) 
      -- CP-element group 480: 	 branch_block_stmt_33/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_677/phi_stmt_677_sources/type_cast_683/SplitProtocol/Sample/$exit
      -- CP-element group 480: 	 branch_block_stmt_33/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_677/phi_stmt_677_sources/type_cast_683/SplitProtocol/Sample/ra
      -- 
    ra_3580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 480_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_683_inst_ack_0, ack => convTranspose_CP_39_elements(480)); -- 
    -- CP-element group 481:  transition  input  bypass 
    -- CP-element group 481: predecessors 
    -- CP-element group 481: 	210 
    -- CP-element group 481: successors 
    -- CP-element group 481: 	482 
    -- CP-element group 481:  members (2) 
      -- CP-element group 481: 	 branch_block_stmt_33/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_677/phi_stmt_677_sources/type_cast_683/SplitProtocol/Update/$exit
      -- CP-element group 481: 	 branch_block_stmt_33/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_677/phi_stmt_677_sources/type_cast_683/SplitProtocol/Update/ca
      -- 
    ca_3585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 481_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_683_inst_ack_1, ack => convTranspose_CP_39_elements(481)); -- 
    -- CP-element group 482:  join  transition  output  bypass 
    -- CP-element group 482: predecessors 
    -- CP-element group 482: 	480 
    -- CP-element group 482: 	481 
    -- CP-element group 482: successors 
    -- CP-element group 482: 	483 
    -- CP-element group 482:  members (6) 
      -- CP-element group 482: 	 branch_block_stmt_33/forx_xbody196_forx_xbody196_PhiReq/$exit
      -- CP-element group 482: 	 branch_block_stmt_33/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_677/$exit
      -- CP-element group 482: 	 branch_block_stmt_33/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_677/phi_stmt_677_sources/$exit
      -- CP-element group 482: 	 branch_block_stmt_33/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_677/phi_stmt_677_sources/type_cast_683/$exit
      -- CP-element group 482: 	 branch_block_stmt_33/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_677/phi_stmt_677_sources/type_cast_683/SplitProtocol/$exit
      -- CP-element group 482: 	 branch_block_stmt_33/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_677/phi_stmt_677_req
      -- 
    phi_stmt_677_req_3586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_677_req_3586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(482), ack => phi_stmt_677_req_1); -- 
    convTranspose_cp_element_group_482: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_482"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(480) & convTranspose_CP_39_elements(481);
      gj_convTranspose_cp_element_group_482 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(482), clk => clk, reset => reset); --
    end block;
    -- CP-element group 483:  merge  transition  place  bypass 
    -- CP-element group 483: predecessors 
    -- CP-element group 483: 	479 
    -- CP-element group 483: 	482 
    -- CP-element group 483: successors 
    -- CP-element group 483: 	484 
    -- CP-element group 483:  members (2) 
      -- CP-element group 483: 	 branch_block_stmt_33/merge_stmt_676_PhiReqMerge
      -- CP-element group 483: 	 branch_block_stmt_33/merge_stmt_676_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(483) <= OrReduce(convTranspose_CP_39_elements(479) & convTranspose_CP_39_elements(482));
    -- CP-element group 484:  fork  transition  place  input  output  bypass 
    -- CP-element group 484: predecessors 
    -- CP-element group 484: 	483 
    -- CP-element group 484: successors 
    -- CP-element group 484: 	180 
    -- CP-element group 484: 	184 
    -- CP-element group 484: 	188 
    -- CP-element group 484: 	192 
    -- CP-element group 484: 	196 
    -- CP-element group 484: 	200 
    -- CP-element group 484: 	204 
    -- CP-element group 484: 	207 
    -- CP-element group 484: 	173 
    -- CP-element group 484: 	176 
    -- CP-element group 484: 	169 
    -- CP-element group 484: 	170 
    -- CP-element group 484: 	172 
    -- CP-element group 484:  members (56) 
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_728_Update/cr
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_728_Update/$entry
      -- CP-element group 484: 	 branch_block_stmt_33/merge_stmt_676__exit__
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839__entry__
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_final_index_sum_regn_Update/req
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_index_scale_1/scale_rename_ack
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_index_scale_1/scale_rename_req
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_final_index_sum_regn_Update/$entry
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_index_scale_1/$exit
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_index_scale_1/$entry
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_710_Update/cr
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_697_Update/cr
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/addr_of_690_complete/req
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_710_Update/$entry
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_697_Update/$entry
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_index_resize_1/index_resize_ack
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/addr_of_690_complete/$entry
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_index_resize_1/index_resize_req
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_final_index_sum_regn_Sample/req
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_index_resize_1/$exit
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_697_update_start_
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_index_resize_1/$entry
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_index_computed_1
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_index_scaled_1
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_final_index_sum_regn_Sample/$entry
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_index_resized_1
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_728_update_start_
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_final_index_sum_regn_update_start
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/addr_of_690_update_start_
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/$entry
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_693_Sample/rr
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_693_Sample/$entry
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_710_update_start_
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_693_sample_start_
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_746_update_start_
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_746_Update/$entry
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_746_Update/cr
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_764_update_start_
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_764_Update/$entry
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_764_Update/cr
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_782_update_start_
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_782_Update/$entry
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_782_Update/cr
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_800_update_start_
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_800_Update/$entry
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_800_Update/cr
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_818_update_start_
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_818_Update/$entry
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_818_Update/cr
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_update_start_
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_Update/$entry
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_Update/word_access_complete/$entry
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_Update/word_access_complete/word_0/$entry
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_Update/word_access_complete/word_0/cr
      -- CP-element group 484: 	 branch_block_stmt_33/merge_stmt_676_PhiAck/$exit
      -- CP-element group 484: 	 branch_block_stmt_33/merge_stmt_676_PhiAck/phi_stmt_677_ack
      -- 
    phi_stmt_677_ack_3591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 484_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_677_ack_0, ack => convTranspose_CP_39_elements(484)); -- 
    cr_1446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(484), ack => type_cast_728_inst_req_1); -- 
    req_1347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(484), ack => array_obj_ref_689_index_offset_req_1); -- 
    cr_1418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(484), ack => type_cast_710_inst_req_1); -- 
    cr_1390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(484), ack => type_cast_697_inst_req_1); -- 
    req_1362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(484), ack => addr_of_690_final_reg_req_1); -- 
    req_1342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(484), ack => array_obj_ref_689_index_offset_req_0); -- 
    rr_1371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(484), ack => RPIPE_ConvTranspose_input_pipe_693_inst_req_0); -- 
    cr_1474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(484), ack => type_cast_746_inst_req_1); -- 
    cr_1502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(484), ack => type_cast_764_inst_req_1); -- 
    cr_1530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(484), ack => type_cast_782_inst_req_1); -- 
    cr_1558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(484), ack => type_cast_800_inst_req_1); -- 
    cr_1586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(484), ack => type_cast_818_inst_req_1); -- 
    cr_1636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(484), ack => ptr_deref_826_store_0_req_1); -- 
    -- CP-element group 485:  merge  fork  transition  place  output  bypass 
    -- CP-element group 485: predecessors 
    -- CP-element group 485: 	209 
    -- CP-element group 485: 	122 
    -- CP-element group 485: successors 
    -- CP-element group 485: 	211 
    -- CP-element group 485: 	212 
    -- CP-element group 485: 	213 
    -- CP-element group 485: 	214 
    -- CP-element group 485: 	215 
    -- CP-element group 485: 	216 
    -- CP-element group 485:  members (25) 
      -- CP-element group 485: 	 branch_block_stmt_33/merge_stmt_848__exit__
      -- CP-element group 485: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876__entry__
      -- CP-element group 485: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/$entry
      -- CP-element group 485: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_851_sample_start_
      -- CP-element group 485: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_851_update_start_
      -- CP-element group 485: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_851_Sample/$entry
      -- CP-element group 485: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_851_Sample/rr
      -- CP-element group 485: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_851_Update/$entry
      -- CP-element group 485: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_851_Update/cr
      -- CP-element group 485: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_855_sample_start_
      -- CP-element group 485: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_855_update_start_
      -- CP-element group 485: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_855_Sample/$entry
      -- CP-element group 485: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_855_Sample/rr
      -- CP-element group 485: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_855_Update/$entry
      -- CP-element group 485: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_855_Update/cr
      -- CP-element group 485: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_859_sample_start_
      -- CP-element group 485: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_859_update_start_
      -- CP-element group 485: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_859_Sample/$entry
      -- CP-element group 485: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_859_Sample/rr
      -- CP-element group 485: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_859_Update/$entry
      -- CP-element group 485: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_859_Update/cr
      -- CP-element group 485: 	 branch_block_stmt_33/merge_stmt_848_PhiReqMerge
      -- CP-element group 485: 	 branch_block_stmt_33/merge_stmt_848_PhiAck/$entry
      -- CP-element group 485: 	 branch_block_stmt_33/merge_stmt_848_PhiAck/$exit
      -- CP-element group 485: 	 branch_block_stmt_33/merge_stmt_848_PhiAck/dummy
      -- 
    rr_1667_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1667_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(485), ack => type_cast_851_inst_req_0); -- 
    cr_1672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(485), ack => type_cast_851_inst_req_1); -- 
    rr_1681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(485), ack => type_cast_855_inst_req_0); -- 
    cr_1686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(485), ack => type_cast_855_inst_req_1); -- 
    rr_1695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(485), ack => type_cast_859_inst_req_0); -- 
    cr_1700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(485), ack => type_cast_859_inst_req_1); -- 
    convTranspose_CP_39_elements(485) <= OrReduce(convTranspose_CP_39_elements(209) & convTranspose_CP_39_elements(122));
    -- CP-element group 486:  transition  output  delay-element  bypass 
    -- CP-element group 486: predecessors 
    -- CP-element group 486: 	221 
    -- CP-element group 486: successors 
    -- CP-element group 486: 	490 
    -- CP-element group 486:  members (5) 
      -- CP-element group 486: 	 branch_block_stmt_33/bbx_xnph508_forx_xbody266_PhiReq/$exit
      -- CP-element group 486: 	 branch_block_stmt_33/bbx_xnph508_forx_xbody266_PhiReq/phi_stmt_921/$exit
      -- CP-element group 486: 	 branch_block_stmt_33/bbx_xnph508_forx_xbody266_PhiReq/phi_stmt_921/phi_stmt_921_sources/$exit
      -- CP-element group 486: 	 branch_block_stmt_33/bbx_xnph508_forx_xbody266_PhiReq/phi_stmt_921/phi_stmt_921_sources/type_cast_927_konst_delay_trans
      -- CP-element group 486: 	 branch_block_stmt_33/bbx_xnph508_forx_xbody266_PhiReq/phi_stmt_921/phi_stmt_921_req
      -- 
    phi_stmt_921_req_3637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_921_req_3637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(486), ack => phi_stmt_921_req_1); -- 
    -- Element group convTranspose_CP_39_elements(486) is a control-delay.
    cp_element_486_delay: control_delay_element  generic map(name => " 486_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(221), ack => convTranspose_CP_39_elements(486), clk => clk, reset =>reset);
    -- CP-element group 487:  transition  input  bypass 
    -- CP-element group 487: predecessors 
    -- CP-element group 487: 	230 
    -- CP-element group 487: successors 
    -- CP-element group 487: 	489 
    -- CP-element group 487:  members (2) 
      -- CP-element group 487: 	 branch_block_stmt_33/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_921/phi_stmt_921_sources/type_cast_924/SplitProtocol/Sample/$exit
      -- CP-element group 487: 	 branch_block_stmt_33/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_921/phi_stmt_921_sources/type_cast_924/SplitProtocol/Sample/ra
      -- 
    ra_3657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 487_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_924_inst_ack_0, ack => convTranspose_CP_39_elements(487)); -- 
    -- CP-element group 488:  transition  input  bypass 
    -- CP-element group 488: predecessors 
    -- CP-element group 488: 	230 
    -- CP-element group 488: successors 
    -- CP-element group 488: 	489 
    -- CP-element group 488:  members (2) 
      -- CP-element group 488: 	 branch_block_stmt_33/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_921/phi_stmt_921_sources/type_cast_924/SplitProtocol/Update/$exit
      -- CP-element group 488: 	 branch_block_stmt_33/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_921/phi_stmt_921_sources/type_cast_924/SplitProtocol/Update/ca
      -- 
    ca_3662_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 488_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_924_inst_ack_1, ack => convTranspose_CP_39_elements(488)); -- 
    -- CP-element group 489:  join  transition  output  bypass 
    -- CP-element group 489: predecessors 
    -- CP-element group 489: 	487 
    -- CP-element group 489: 	488 
    -- CP-element group 489: successors 
    -- CP-element group 489: 	490 
    -- CP-element group 489:  members (6) 
      -- CP-element group 489: 	 branch_block_stmt_33/forx_xbody266_forx_xbody266_PhiReq/$exit
      -- CP-element group 489: 	 branch_block_stmt_33/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_921/$exit
      -- CP-element group 489: 	 branch_block_stmt_33/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_921/phi_stmt_921_sources/$exit
      -- CP-element group 489: 	 branch_block_stmt_33/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_921/phi_stmt_921_sources/type_cast_924/$exit
      -- CP-element group 489: 	 branch_block_stmt_33/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_921/phi_stmt_921_sources/type_cast_924/SplitProtocol/$exit
      -- CP-element group 489: 	 branch_block_stmt_33/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_921/phi_stmt_921_req
      -- 
    phi_stmt_921_req_3663_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_921_req_3663_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(489), ack => phi_stmt_921_req_0); -- 
    convTranspose_cp_element_group_489: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_489"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(487) & convTranspose_CP_39_elements(488);
      gj_convTranspose_cp_element_group_489 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(489), clk => clk, reset => reset); --
    end block;
    -- CP-element group 490:  merge  transition  place  bypass 
    -- CP-element group 490: predecessors 
    -- CP-element group 490: 	486 
    -- CP-element group 490: 	489 
    -- CP-element group 490: successors 
    -- CP-element group 490: 	491 
    -- CP-element group 490:  members (2) 
      -- CP-element group 490: 	 branch_block_stmt_33/merge_stmt_920_PhiReqMerge
      -- CP-element group 490: 	 branch_block_stmt_33/merge_stmt_920_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(490) <= OrReduce(convTranspose_CP_39_elements(486) & convTranspose_CP_39_elements(489));
    -- CP-element group 491:  fork  transition  place  input  output  bypass 
    -- CP-element group 491: predecessors 
    -- CP-element group 491: 	490 
    -- CP-element group 491: successors 
    -- CP-element group 491: 	222 
    -- CP-element group 491: 	223 
    -- CP-element group 491: 	225 
    -- CP-element group 491: 	227 
    -- CP-element group 491:  members (29) 
      -- CP-element group 491: 	 branch_block_stmt_33/merge_stmt_920__exit__
      -- CP-element group 491: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951__entry__
      -- CP-element group 491: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/$entry
      -- CP-element group 491: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/addr_of_934_update_start_
      -- CP-element group 491: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_index_resized_1
      -- CP-element group 491: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_index_scaled_1
      -- CP-element group 491: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_index_computed_1
      -- CP-element group 491: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_index_resize_1/$entry
      -- CP-element group 491: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_index_resize_1/$exit
      -- CP-element group 491: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_index_resize_1/index_resize_req
      -- CP-element group 491: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_index_resize_1/index_resize_ack
      -- CP-element group 491: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_index_scale_1/$entry
      -- CP-element group 491: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_index_scale_1/$exit
      -- CP-element group 491: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_index_scale_1/scale_rename_req
      -- CP-element group 491: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_index_scale_1/scale_rename_ack
      -- CP-element group 491: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_final_index_sum_regn_update_start
      -- CP-element group 491: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_final_index_sum_regn_Sample/$entry
      -- CP-element group 491: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_final_index_sum_regn_Sample/req
      -- CP-element group 491: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_final_index_sum_regn_Update/$entry
      -- CP-element group 491: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_final_index_sum_regn_Update/req
      -- CP-element group 491: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/addr_of_934_complete/$entry
      -- CP-element group 491: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/addr_of_934_complete/req
      -- CP-element group 491: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_update_start_
      -- CP-element group 491: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_Update/$entry
      -- CP-element group 491: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_Update/word_access_complete/$entry
      -- CP-element group 491: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_Update/word_access_complete/word_0/$entry
      -- CP-element group 491: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_Update/word_access_complete/word_0/cr
      -- CP-element group 491: 	 branch_block_stmt_33/merge_stmt_920_PhiAck/$exit
      -- CP-element group 491: 	 branch_block_stmt_33/merge_stmt_920_PhiAck/phi_stmt_921_ack
      -- 
    phi_stmt_921_ack_3668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 491_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_921_ack_0, ack => convTranspose_CP_39_elements(491)); -- 
    req_1765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(491), ack => array_obj_ref_933_index_offset_req_0); -- 
    req_1770_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1770_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(491), ack => array_obj_ref_933_index_offset_req_1); -- 
    req_1785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(491), ack => addr_of_934_final_reg_req_1); -- 
    cr_1835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(491), ack => ptr_deref_937_store_0_req_1); -- 
    -- CP-element group 492:  merge  fork  transition  place  output  bypass 
    -- CP-element group 492: predecessors 
    -- CP-element group 492: 	219 
    -- CP-element group 492: 	229 
    -- CP-element group 492: successors 
    -- CP-element group 492: 	231 
    -- CP-element group 492: 	232 
    -- CP-element group 492: 	234 
    -- CP-element group 492:  members (16) 
      -- CP-element group 492: 	 branch_block_stmt_33/merge_stmt_960__exit__
      -- CP-element group 492: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_969__entry__
      -- CP-element group 492: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_969/$entry
      -- CP-element group 492: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_969/call_stmt_963_sample_start_
      -- CP-element group 492: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_969/call_stmt_963_update_start_
      -- CP-element group 492: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_969/call_stmt_963_Sample/$entry
      -- CP-element group 492: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_969/call_stmt_963_Sample/crr
      -- CP-element group 492: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_969/call_stmt_963_Update/$entry
      -- CP-element group 492: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_969/call_stmt_963_Update/ccr
      -- CP-element group 492: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_969/type_cast_968_update_start_
      -- CP-element group 492: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_969/type_cast_968_Update/$entry
      -- CP-element group 492: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_969/type_cast_968_Update/cr
      -- CP-element group 492: 	 branch_block_stmt_33/merge_stmt_960_PhiReqMerge
      -- CP-element group 492: 	 branch_block_stmt_33/merge_stmt_960_PhiAck/$entry
      -- CP-element group 492: 	 branch_block_stmt_33/merge_stmt_960_PhiAck/$exit
      -- CP-element group 492: 	 branch_block_stmt_33/merge_stmt_960_PhiAck/dummy
      -- 
    crr_1866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(492), ack => call_stmt_963_call_req_0); -- 
    ccr_1871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(492), ack => call_stmt_963_call_req_1); -- 
    cr_1885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(492), ack => type_cast_968_inst_req_1); -- 
    convTranspose_CP_39_elements(492) <= OrReduce(convTranspose_CP_39_elements(219) & convTranspose_CP_39_elements(229));
    -- CP-element group 493:  transition  output  delay-element  bypass 
    -- CP-element group 493: predecessors 
    -- CP-element group 493: 	423 
    -- CP-element group 493: successors 
    -- CP-element group 493: 	497 
    -- CP-element group 493:  members (5) 
      -- CP-element group 493: 	 branch_block_stmt_33/bbx_xnph_forx_xbody428_PhiReq/$exit
      -- CP-element group 493: 	 branch_block_stmt_33/bbx_xnph_forx_xbody428_PhiReq/phi_stmt_1354/$exit
      -- CP-element group 493: 	 branch_block_stmt_33/bbx_xnph_forx_xbody428_PhiReq/phi_stmt_1354/phi_stmt_1354_sources/$exit
      -- CP-element group 493: 	 branch_block_stmt_33/bbx_xnph_forx_xbody428_PhiReq/phi_stmt_1354/phi_stmt_1354_sources/type_cast_1358_konst_delay_trans
      -- CP-element group 493: 	 branch_block_stmt_33/bbx_xnph_forx_xbody428_PhiReq/phi_stmt_1354/phi_stmt_1354_req
      -- 
    phi_stmt_1354_req_3714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1354_req_3714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(493), ack => phi_stmt_1354_req_0); -- 
    -- Element group convTranspose_CP_39_elements(493) is a control-delay.
    cp_element_493_delay: control_delay_element  generic map(name => " 493_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(423), ack => convTranspose_CP_39_elements(493), clk => clk, reset =>reset);
    -- CP-element group 494:  transition  input  bypass 
    -- CP-element group 494: predecessors 
    -- CP-element group 494: 	471 
    -- CP-element group 494: successors 
    -- CP-element group 494: 	496 
    -- CP-element group 494:  members (2) 
      -- CP-element group 494: 	 branch_block_stmt_33/forx_xbody428_forx_xbody428_PhiReq/phi_stmt_1354/phi_stmt_1354_sources/type_cast_1360/SplitProtocol/Sample/$exit
      -- CP-element group 494: 	 branch_block_stmt_33/forx_xbody428_forx_xbody428_PhiReq/phi_stmt_1354/phi_stmt_1354_sources/type_cast_1360/SplitProtocol/Sample/ra
      -- 
    ra_3734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 494_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1360_inst_ack_0, ack => convTranspose_CP_39_elements(494)); -- 
    -- CP-element group 495:  transition  input  bypass 
    -- CP-element group 495: predecessors 
    -- CP-element group 495: 	471 
    -- CP-element group 495: successors 
    -- CP-element group 495: 	496 
    -- CP-element group 495:  members (2) 
      -- CP-element group 495: 	 branch_block_stmt_33/forx_xbody428_forx_xbody428_PhiReq/phi_stmt_1354/phi_stmt_1354_sources/type_cast_1360/SplitProtocol/Update/$exit
      -- CP-element group 495: 	 branch_block_stmt_33/forx_xbody428_forx_xbody428_PhiReq/phi_stmt_1354/phi_stmt_1354_sources/type_cast_1360/SplitProtocol/Update/ca
      -- 
    ca_3739_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 495_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1360_inst_ack_1, ack => convTranspose_CP_39_elements(495)); -- 
    -- CP-element group 496:  join  transition  output  bypass 
    -- CP-element group 496: predecessors 
    -- CP-element group 496: 	494 
    -- CP-element group 496: 	495 
    -- CP-element group 496: successors 
    -- CP-element group 496: 	497 
    -- CP-element group 496:  members (6) 
      -- CP-element group 496: 	 branch_block_stmt_33/forx_xbody428_forx_xbody428_PhiReq/$exit
      -- CP-element group 496: 	 branch_block_stmt_33/forx_xbody428_forx_xbody428_PhiReq/phi_stmt_1354/$exit
      -- CP-element group 496: 	 branch_block_stmt_33/forx_xbody428_forx_xbody428_PhiReq/phi_stmt_1354/phi_stmt_1354_sources/$exit
      -- CP-element group 496: 	 branch_block_stmt_33/forx_xbody428_forx_xbody428_PhiReq/phi_stmt_1354/phi_stmt_1354_sources/type_cast_1360/$exit
      -- CP-element group 496: 	 branch_block_stmt_33/forx_xbody428_forx_xbody428_PhiReq/phi_stmt_1354/phi_stmt_1354_sources/type_cast_1360/SplitProtocol/$exit
      -- CP-element group 496: 	 branch_block_stmt_33/forx_xbody428_forx_xbody428_PhiReq/phi_stmt_1354/phi_stmt_1354_req
      -- 
    phi_stmt_1354_req_3740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1354_req_3740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(496), ack => phi_stmt_1354_req_1); -- 
    convTranspose_cp_element_group_496: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_496"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(494) & convTranspose_CP_39_elements(495);
      gj_convTranspose_cp_element_group_496 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(496), clk => clk, reset => reset); --
    end block;
    -- CP-element group 497:  merge  transition  place  bypass 
    -- CP-element group 497: predecessors 
    -- CP-element group 497: 	493 
    -- CP-element group 497: 	496 
    -- CP-element group 497: successors 
    -- CP-element group 497: 	498 
    -- CP-element group 497:  members (2) 
      -- CP-element group 497: 	 branch_block_stmt_33/merge_stmt_1353_PhiReqMerge
      -- CP-element group 497: 	 branch_block_stmt_33/merge_stmt_1353_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(497) <= OrReduce(convTranspose_CP_39_elements(493) & convTranspose_CP_39_elements(496));
    -- CP-element group 498:  fork  transition  place  input  output  bypass 
    -- CP-element group 498: predecessors 
    -- CP-element group 498: 	497 
    -- CP-element group 498: successors 
    -- CP-element group 498: 	424 
    -- CP-element group 498: 	425 
    -- CP-element group 498: 	427 
    -- CP-element group 498: 	429 
    -- CP-element group 498: 	431 
    -- CP-element group 498: 	433 
    -- CP-element group 498: 	435 
    -- CP-element group 498: 	437 
    -- CP-element group 498: 	439 
    -- CP-element group 498: 	441 
    -- CP-element group 498: 	443 
    -- CP-element group 498: 	445 
    -- CP-element group 498:  members (53) 
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1425_Update/$entry
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/array_obj_ref_1366_index_resize_1/$entry
      -- CP-element group 498: 	 branch_block_stmt_33/merge_stmt_1353__exit__
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481__entry__
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1445_update_start_
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1395_Update/cr
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/array_obj_ref_1366_index_scale_1/$exit
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/array_obj_ref_1366_index_computed_1
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1425_update_start_
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1375_Update/$entry
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1425_Update/cr
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1405_update_start_
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/array_obj_ref_1366_index_scaled_1
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/array_obj_ref_1366_index_scale_1/$entry
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/array_obj_ref_1366_index_resize_1/$exit
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1395_Update/$entry
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/array_obj_ref_1366_index_resize_1/index_resize_req
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/array_obj_ref_1366_index_resized_1
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/array_obj_ref_1366_index_resize_1/index_resize_ack
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/addr_of_1367_complete/$entry
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/array_obj_ref_1366_index_scale_1/scale_rename_req
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1375_Update/cr
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/array_obj_ref_1366_index_scale_1/scale_rename_ack
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/array_obj_ref_1366_final_index_sum_regn_update_start
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/array_obj_ref_1366_final_index_sum_regn_Sample/$entry
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/array_obj_ref_1366_final_index_sum_regn_Sample/req
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/array_obj_ref_1366_final_index_sum_regn_Update/$entry
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/array_obj_ref_1366_final_index_sum_regn_Update/req
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/addr_of_1367_complete/req
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1405_Update/$entry
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1435_update_start_
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1375_update_start_
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1395_update_start_
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/addr_of_1367_update_start_
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1435_Update/cr
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/$entry
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1385_Update/cr
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1385_Update/$entry
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/ptr_deref_1371_Update/word_access_complete/word_0/cr
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/ptr_deref_1371_Update/word_access_complete/word_0/$entry
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1415_Update/cr
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/ptr_deref_1371_Update/word_access_complete/$entry
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/ptr_deref_1371_Update/$entry
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1415_Update/$entry
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1435_Update/$entry
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1415_update_start_
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1385_update_start_
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1445_Update/cr
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1405_Update/cr
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/ptr_deref_1371_update_start_
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1368_to_assign_stmt_1481/type_cast_1445_Update/$entry
      -- CP-element group 498: 	 branch_block_stmt_33/merge_stmt_1353_PhiAck/$exit
      -- CP-element group 498: 	 branch_block_stmt_33/merge_stmt_1353_PhiAck/phi_stmt_1354_ack
      -- 
    phi_stmt_1354_ack_3745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 498_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1354_ack_0, ack => convTranspose_CP_39_elements(498)); -- 
    cr_3258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(498), ack => type_cast_1395_inst_req_1); -- 
    cr_3300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(498), ack => type_cast_1425_inst_req_1); -- 
    cr_3230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(498), ack => type_cast_1375_inst_req_1); -- 
    req_3146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(498), ack => array_obj_ref_1366_index_offset_req_0); -- 
    req_3151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(498), ack => array_obj_ref_1366_index_offset_req_1); -- 
    req_3166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(498), ack => addr_of_1367_final_reg_req_1); -- 
    cr_3314_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3314_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(498), ack => type_cast_1435_inst_req_1); -- 
    cr_3244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(498), ack => type_cast_1385_inst_req_1); -- 
    cr_3211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(498), ack => ptr_deref_1371_load_0_req_1); -- 
    cr_3286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(498), ack => type_cast_1415_inst_req_1); -- 
    cr_3328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(498), ack => type_cast_1445_inst_req_1); -- 
    cr_3272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(498), ack => type_cast_1405_inst_req_1); -- 
    -- CP-element group 499:  merge  transition  place  bypass 
    -- CP-element group 499: predecessors 
    -- CP-element group 499: 	421 
    -- CP-element group 499: 	470 
    -- CP-element group 499: successors 
    -- CP-element group 499:  members (16) 
      -- CP-element group 499: 	 $exit
      -- CP-element group 499: 	 branch_block_stmt_33/$exit
      -- CP-element group 499: 	 branch_block_stmt_33/branch_block_stmt_33__exit__
      -- CP-element group 499: 	 branch_block_stmt_33/merge_stmt_1490__exit__
      -- CP-element group 499: 	 branch_block_stmt_33/return__
      -- CP-element group 499: 	 branch_block_stmt_33/merge_stmt_1492__exit__
      -- CP-element group 499: 	 branch_block_stmt_33/merge_stmt_1490_PhiReqMerge
      -- CP-element group 499: 	 branch_block_stmt_33/merge_stmt_1490_PhiAck/$entry
      -- CP-element group 499: 	 branch_block_stmt_33/merge_stmt_1490_PhiAck/$exit
      -- CP-element group 499: 	 branch_block_stmt_33/merge_stmt_1490_PhiAck/dummy
      -- CP-element group 499: 	 branch_block_stmt_33/return___PhiReq/$entry
      -- CP-element group 499: 	 branch_block_stmt_33/return___PhiReq/$exit
      -- CP-element group 499: 	 branch_block_stmt_33/merge_stmt_1492_PhiReqMerge
      -- CP-element group 499: 	 branch_block_stmt_33/merge_stmt_1492_PhiAck/$entry
      -- CP-element group 499: 	 branch_block_stmt_33/merge_stmt_1492_PhiAck/$exit
      -- CP-element group 499: 	 branch_block_stmt_33/merge_stmt_1492_PhiAck/dummy
      -- 
    convTranspose_CP_39_elements(499) <= OrReduce(convTranspose_CP_39_elements(421) & convTranspose_CP_39_elements(470));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar526_932_resized : std_logic_vector(13 downto 0);
    signal R_indvar526_932_scaled : std_logic_vector(13 downto 0);
    signal R_indvar540_688_resized : std_logic_vector(10 downto 0);
    signal R_indvar540_688_scaled : std_logic_vector(10 downto 0);
    signal R_indvar556_481_resized : std_logic_vector(13 downto 0);
    signal R_indvar556_481_scaled : std_logic_vector(13 downto 0);
    signal R_indvar_1365_resized : std_logic_vector(13 downto 0);
    signal R_indvar_1365_scaled : std_logic_vector(13 downto 0);
    signal add108_334 : std_logic_vector(15 downto 0);
    signal add117_359 : std_logic_vector(15 downto 0);
    signal add126_384 : std_logic_vector(15 downto 0);
    signal add12_83 : std_logic_vector(15 downto 0);
    signal add135_409 : std_logic_vector(15 downto 0);
    signal add150_509 : std_logic_vector(63 downto 0);
    signal add156_527 : std_logic_vector(63 downto 0);
    signal add162_545 : std_logic_vector(63 downto 0);
    signal add168_563 : std_logic_vector(63 downto 0);
    signal add174_581 : std_logic_vector(63 downto 0);
    signal add180_599 : std_logic_vector(63 downto 0);
    signal add186_617 : std_logic_vector(63 downto 0);
    signal add206_716 : std_logic_vector(63 downto 0);
    signal add212_734 : std_logic_vector(63 downto 0);
    signal add218_752 : std_logic_vector(63 downto 0);
    signal add21_108 : std_logic_vector(15 downto 0);
    signal add224_770 : std_logic_vector(63 downto 0);
    signal add230_788 : std_logic_vector(63 downto 0);
    signal add236_806 : std_logic_vector(63 downto 0);
    signal add242_824 : std_logic_vector(63 downto 0);
    signal add30_133 : std_logic_vector(15 downto 0);
    signal add39_158 : std_logic_vector(15 downto 0);
    signal add48_183 : std_logic_vector(15 downto 0);
    signal add57_208 : std_logic_vector(15 downto 0);
    signal add74_248 : std_logic_vector(31 downto 0);
    signal add79_253 : std_logic_vector(31 downto 0);
    signal add99_309 : std_logic_vector(15 downto 0);
    signal add_58 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1366_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1366_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1366_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1366_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1366_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1366_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_482_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_482_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_482_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_482_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_482_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_482_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_689_constant_part_of_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_689_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_689_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_689_offset_scale_factor_1 : std_logic_vector(10 downto 0);
    signal array_obj_ref_689_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_689_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_933_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_933_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_933_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_933_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_933_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_933_root_address : std_logic_vector(13 downto 0);
    signal arrayidx246_691 : std_logic_vector(31 downto 0);
    signal arrayidx269_935 : std_logic_vector(31 downto 0);
    signal arrayidx433_1368 : std_logic_vector(31 downto 0);
    signal arrayidx_484 : std_logic_vector(31 downto 0);
    signal call101_312 : std_logic_vector(7 downto 0);
    signal call106_325 : std_logic_vector(7 downto 0);
    signal call10_74 : std_logic_vector(7 downto 0);
    signal call110_337 : std_logic_vector(7 downto 0);
    signal call115_350 : std_logic_vector(7 downto 0);
    signal call119_362 : std_logic_vector(7 downto 0);
    signal call124_375 : std_logic_vector(7 downto 0);
    signal call128_387 : std_logic_vector(7 downto 0);
    signal call133_400 : std_logic_vector(7 downto 0);
    signal call143_487 : std_logic_vector(7 downto 0);
    signal call147_500 : std_logic_vector(7 downto 0);
    signal call14_86 : std_logic_vector(7 downto 0);
    signal call153_518 : std_logic_vector(7 downto 0);
    signal call159_536 : std_logic_vector(7 downto 0);
    signal call165_554 : std_logic_vector(7 downto 0);
    signal call171_572 : std_logic_vector(7 downto 0);
    signal call177_590 : std_logic_vector(7 downto 0);
    signal call183_608 : std_logic_vector(7 downto 0);
    signal call199_694 : std_logic_vector(7 downto 0);
    signal call19_99 : std_logic_vector(7 downto 0);
    signal call203_707 : std_logic_vector(7 downto 0);
    signal call209_725 : std_logic_vector(7 downto 0);
    signal call215_743 : std_logic_vector(7 downto 0);
    signal call221_761 : std_logic_vector(7 downto 0);
    signal call227_779 : std_logic_vector(7 downto 0);
    signal call233_797 : std_logic_vector(7 downto 0);
    signal call239_815 : std_logic_vector(7 downto 0);
    signal call23_111 : std_logic_vector(7 downto 0);
    signal call275_963 : std_logic_vector(63 downto 0);
    signal call28_124 : std_logic_vector(7 downto 0);
    signal call2_49 : std_logic_vector(7 downto 0);
    signal call32_136 : std_logic_vector(7 downto 0);
    signal call346_1185 : std_logic_vector(15 downto 0);
    signal call348_1188 : std_logic_vector(15 downto 0);
    signal call350_1191 : std_logic_vector(15 downto 0);
    signal call352_1194 : std_logic_vector(15 downto 0);
    signal call354_1197 : std_logic_vector(63 downto 0);
    signal call37_149 : std_logic_vector(7 downto 0);
    signal call41_161 : std_logic_vector(7 downto 0);
    signal call46_174 : std_logic_vector(7 downto 0);
    signal call50_186 : std_logic_vector(7 downto 0);
    signal call55_199 : std_logic_vector(7 downto 0);
    signal call5_61 : std_logic_vector(7 downto 0);
    signal call92_287 : std_logic_vector(7 downto 0);
    signal call97_300 : std_logic_vector(7 downto 0);
    signal call_36 : std_logic_vector(7 downto 0);
    signal cmp194510_431 : std_logic_vector(0 downto 0);
    signal cmp264506_876 : std_logic_vector(0 downto 0);
    signal cmp514_416 : std_logic_vector(0 downto 0);
    signal conv104_316 : std_logic_vector(15 downto 0);
    signal conv107_329 : std_logic_vector(15 downto 0);
    signal conv113_341 : std_logic_vector(15 downto 0);
    signal conv116_354 : std_logic_vector(15 downto 0);
    signal conv11_78 : std_logic_vector(15 downto 0);
    signal conv122_366 : std_logic_vector(15 downto 0);
    signal conv125_379 : std_logic_vector(15 downto 0);
    signal conv131_391 : std_logic_vector(15 downto 0);
    signal conv134_404 : std_logic_vector(15 downto 0);
    signal conv144_491 : std_logic_vector(63 downto 0);
    signal conv149_504 : std_logic_vector(63 downto 0);
    signal conv155_522 : std_logic_vector(63 downto 0);
    signal conv161_540 : std_logic_vector(63 downto 0);
    signal conv167_558 : std_logic_vector(63 downto 0);
    signal conv173_576 : std_logic_vector(63 downto 0);
    signal conv179_594 : std_logic_vector(63 downto 0);
    signal conv17_90 : std_logic_vector(15 downto 0);
    signal conv185_612 : std_logic_vector(63 downto 0);
    signal conv1_40 : std_logic_vector(15 downto 0);
    signal conv200_698 : std_logic_vector(63 downto 0);
    signal conv205_711 : std_logic_vector(63 downto 0);
    signal conv20_103 : std_logic_vector(15 downto 0);
    signal conv211_729 : std_logic_vector(63 downto 0);
    signal conv217_747 : std_logic_vector(63 downto 0);
    signal conv223_765 : std_logic_vector(63 downto 0);
    signal conv229_783 : std_logic_vector(63 downto 0);
    signal conv235_801 : std_logic_vector(63 downto 0);
    signal conv241_819 : std_logic_vector(63 downto 0);
    signal conv253_852 : std_logic_vector(31 downto 0);
    signal conv255_856 : std_logic_vector(31 downto 0);
    signal conv258_860 : std_logic_vector(31 downto 0);
    signal conv26_115 : std_logic_vector(15 downto 0);
    signal conv276_969 : std_logic_vector(63 downto 0);
    signal conv29_128 : std_logic_vector(15 downto 0);
    signal conv305_1051 : std_logic_vector(15 downto 0);
    signal conv307_1058 : std_logic_vector(15 downto 0);
    signal conv322_1107 : std_logic_vector(15 downto 0);
    signal conv324_1114 : std_logic_vector(15 downto 0);
    signal conv339_1163 : std_logic_vector(15 downto 0);
    signal conv341_1170 : std_logic_vector(15 downto 0);
    signal conv355_1202 : std_logic_vector(63 downto 0);
    signal conv35_140 : std_logic_vector(15 downto 0);
    signal conv362_1214 : std_logic_vector(7 downto 0);
    signal conv368_1224 : std_logic_vector(7 downto 0);
    signal conv374_1234 : std_logic_vector(7 downto 0);
    signal conv380_1244 : std_logic_vector(7 downto 0);
    signal conv386_1254 : std_logic_vector(7 downto 0);
    signal conv38_153 : std_logic_vector(15 downto 0);
    signal conv392_1264 : std_logic_vector(7 downto 0);
    signal conv398_1274 : std_logic_vector(7 downto 0);
    signal conv3_53 : std_logic_vector(15 downto 0);
    signal conv404_1284 : std_logic_vector(7 downto 0);
    signal conv438_1376 : std_logic_vector(7 downto 0);
    signal conv444_1386 : std_logic_vector(7 downto 0);
    signal conv44_165 : std_logic_vector(15 downto 0);
    signal conv450_1396 : std_logic_vector(7 downto 0);
    signal conv456_1406 : std_logic_vector(7 downto 0);
    signal conv462_1416 : std_logic_vector(7 downto 0);
    signal conv468_1426 : std_logic_vector(7 downto 0);
    signal conv474_1436 : std_logic_vector(7 downto 0);
    signal conv47_178 : std_logic_vector(15 downto 0);
    signal conv480_1446 : std_logic_vector(7 downto 0);
    signal conv53_190 : std_logic_vector(15 downto 0);
    signal conv56_203 : std_logic_vector(15 downto 0);
    signal conv61_212 : std_logic_vector(31 downto 0);
    signal conv63_216 : std_logic_vector(31 downto 0);
    signal conv65_220 : std_logic_vector(31 downto 0);
    signal conv82_257 : std_logic_vector(31 downto 0);
    signal conv84_261 : std_logic_vector(31 downto 0);
    signal conv87_265 : std_logic_vector(31 downto 0);
    signal conv8_65 : std_logic_vector(15 downto 0);
    signal conv90_269 : std_logic_vector(31 downto 0);
    signal conv95_291 : std_logic_vector(15 downto 0);
    signal conv98_304 : std_logic_vector(15 downto 0);
    signal exitcond1_1481 : std_logic_vector(0 downto 0);
    signal exitcond2_839 : std_logic_vector(0 downto 0);
    signal exitcond3_632 : std_logic_vector(0 downto 0);
    signal exitcond_951 : std_logic_vector(0 downto 0);
    signal iNsTr_14_242 : std_logic_vector(31 downto 0);
    signal iNsTr_197_1338 : std_logic_vector(63 downto 0);
    signal iNsTr_26_454 : std_logic_vector(63 downto 0);
    signal iNsTr_39_661 : std_logic_vector(63 downto 0);
    signal iNsTr_53_905 : std_logic_vector(63 downto 0);
    signal indvar526_921 : std_logic_vector(63 downto 0);
    signal indvar540_677 : std_logic_vector(63 downto 0);
    signal indvar556_470 : std_logic_vector(63 downto 0);
    signal indvar_1354 : std_logic_vector(63 downto 0);
    signal indvarx_xnext527_946 : std_logic_vector(63 downto 0);
    signal indvarx_xnext541_834 : std_logic_vector(63 downto 0);
    signal indvarx_xnext557_627 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1476 : std_logic_vector(63 downto 0);
    signal mul256_865 : std_logic_vector(31 downto 0);
    signal mul259_870 : std_logic_vector(31 downto 0);
    signal mul66_230 : std_logic_vector(31 downto 0);
    signal mul85_274 : std_logic_vector(31 downto 0);
    signal mul88_279 : std_logic_vector(31 downto 0);
    signal mul91_284 : std_logic_vector(31 downto 0);
    signal mul_225 : std_logic_vector(31 downto 0);
    signal ptr_deref_1371_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1371_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1371_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1371_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1371_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_619_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_619_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_619_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_619_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_619_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_619_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_826_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_826_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_826_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_826_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_826_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_826_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_937_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_937_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_937_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_937_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_937_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_937_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl105_322 : std_logic_vector(15 downto 0);
    signal shl114_347 : std_logic_vector(15 downto 0);
    signal shl123_372 : std_logic_vector(15 downto 0);
    signal shl132_397 : std_logic_vector(15 downto 0);
    signal shl146_497 : std_logic_vector(63 downto 0);
    signal shl152_515 : std_logic_vector(63 downto 0);
    signal shl158_533 : std_logic_vector(63 downto 0);
    signal shl164_551 : std_logic_vector(63 downto 0);
    signal shl170_569 : std_logic_vector(63 downto 0);
    signal shl176_587 : std_logic_vector(63 downto 0);
    signal shl182_605 : std_logic_vector(63 downto 0);
    signal shl18_96 : std_logic_vector(15 downto 0);
    signal shl202_704 : std_logic_vector(63 downto 0);
    signal shl208_722 : std_logic_vector(63 downto 0);
    signal shl214_740 : std_logic_vector(63 downto 0);
    signal shl220_758 : std_logic_vector(63 downto 0);
    signal shl226_776 : std_logic_vector(63 downto 0);
    signal shl232_794 : std_logic_vector(63 downto 0);
    signal shl238_812 : std_logic_vector(63 downto 0);
    signal shl27_121 : std_logic_vector(15 downto 0);
    signal shl36_146 : std_logic_vector(15 downto 0);
    signal shl45_171 : std_logic_vector(15 downto 0);
    signal shl54_196 : std_logic_vector(15 downto 0);
    signal shl96_297 : std_logic_vector(15 downto 0);
    signal shl9_71 : std_logic_vector(15 downto 0);
    signal shl_46 : std_logic_vector(15 downto 0);
    signal shr304_1047 : std_logic_vector(31 downto 0);
    signal shr321_1103 : std_logic_vector(31 downto 0);
    signal shr338_1159 : std_logic_vector(31 downto 0);
    signal shr365_1220 : std_logic_vector(63 downto 0);
    signal shr371_1230 : std_logic_vector(63 downto 0);
    signal shr377_1240 : std_logic_vector(63 downto 0);
    signal shr383_1250 : std_logic_vector(63 downto 0);
    signal shr389_1260 : std_logic_vector(63 downto 0);
    signal shr395_1270 : std_logic_vector(63 downto 0);
    signal shr401_1280 : std_logic_vector(63 downto 0);
    signal shr441_1382 : std_logic_vector(63 downto 0);
    signal shr447_1392 : std_logic_vector(63 downto 0);
    signal shr453_1402 : std_logic_vector(63 downto 0);
    signal shr459_1412 : std_logic_vector(63 downto 0);
    signal shr465_1422 : std_logic_vector(63 downto 0);
    signal shr471_1432 : std_logic_vector(63 downto 0);
    signal shr477_1442 : std_logic_vector(63 downto 0);
    signal shr_236 : std_logic_vector(31 downto 0);
    signal sub_1207 : std_logic_vector(63 downto 0);
    signal tmp434_1372 : std_logic_vector(63 downto 0);
    signal tmp521_1322 : std_logic_vector(31 downto 0);
    signal tmp521x_xop_1334 : std_logic_vector(31 downto 0);
    signal tmp522_1328 : std_logic_vector(0 downto 0);
    signal tmp525_1351 : std_logic_vector(63 downto 0);
    signal tmp533_889 : std_logic_vector(31 downto 0);
    signal tmp533x_xop_901 : std_logic_vector(31 downto 0);
    signal tmp534_895 : std_logic_vector(0 downto 0);
    signal tmp538_918 : std_logic_vector(63 downto 0);
    signal tmp549_645 : std_logic_vector(31 downto 0);
    signal tmp549x_xop_657 : std_logic_vector(31 downto 0);
    signal tmp550_651 : std_logic_vector(0 downto 0);
    signal tmp554_674 : std_logic_vector(63 downto 0);
    signal tmp563x_xop_450 : std_logic_vector(31 downto 0);
    signal tmp564_444 : std_logic_vector(0 downto 0);
    signal tmp568_467 : std_logic_vector(63 downto 0);
    signal type_cast_1000_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1004_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1045_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1101_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1157_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_119_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1200_wire : std_logic_vector(63 downto 0);
    signal type_cast_1218_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1228_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1238_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1248_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1258_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1268_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1278_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1320_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1326_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1332_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1342_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1349_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1358_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1360_wire : std_logic_vector(63 downto 0);
    signal type_cast_1380_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1390_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1400_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1410_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1420_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1430_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1440_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_144_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1474_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_169_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_194_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_234_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_240_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_246_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_295_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_320_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_345_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_370_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_395_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_413_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_429_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_442_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_448_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_44_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_458_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_465_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_474_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_476_wire : std_logic_vector(63 downto 0);
    signal type_cast_495_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_513_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_531_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_549_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_567_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_585_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_603_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_625_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_643_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_649_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_655_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_665_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_672_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_681_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_683_wire : std_logic_vector(63 downto 0);
    signal type_cast_69_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_702_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_720_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_738_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_756_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_774_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_792_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_810_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_832_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_874_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_887_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_893_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_899_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_909_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_916_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_924_wire : std_logic_vector(63 downto 0);
    signal type_cast_927_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_939_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_944_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_94_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_967_wire : std_logic_vector(63 downto 0);
    signal xx_xop570_911 : std_logic_vector(63 downto 0);
    signal xx_xop571_667 : std_logic_vector(63 downto 0);
    signal xx_xop572_460 : std_logic_vector(63 downto 0);
    signal xx_xop_1344 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1366_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1366_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1366_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1366_resized_base_address <= "00000000000000";
    array_obj_ref_482_constant_part_of_offset <= "00000000000000";
    array_obj_ref_482_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_482_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_482_resized_base_address <= "00000000000000";
    array_obj_ref_689_constant_part_of_offset <= "00000100010";
    array_obj_ref_689_offset_scale_factor_0 <= "10000000000";
    array_obj_ref_689_offset_scale_factor_1 <= "00000000001";
    array_obj_ref_689_resized_base_address <= "00000000000";
    array_obj_ref_933_constant_part_of_offset <= "00000000000000";
    array_obj_ref_933_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_933_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_933_resized_base_address <= "00000000000000";
    ptr_deref_1371_word_offset_0 <= "00000000000000";
    ptr_deref_619_word_offset_0 <= "00000000000000";
    ptr_deref_826_word_offset_0 <= "00000000000";
    ptr_deref_937_word_offset_0 <= "00000000000000";
    type_cast_1000_wire_constant <= "0000000000000000";
    type_cast_1004_wire_constant <= "0000000000000000";
    type_cast_1045_wire_constant <= "00000000000000000000000000010010";
    type_cast_1101_wire_constant <= "00000000000000000000000000010001";
    type_cast_1157_wire_constant <= "00000000000000000000000000010000";
    type_cast_119_wire_constant <= "0000000000001000";
    type_cast_1218_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1228_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1238_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1248_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1258_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1268_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1278_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1320_wire_constant <= "00000000000000000000000000000010";
    type_cast_1326_wire_constant <= "00000000000000000000000000000001";
    type_cast_1332_wire_constant <= "11111111111111111111111111111111";
    type_cast_1342_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1349_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1358_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1380_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1390_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1400_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1410_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1420_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1430_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1440_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_144_wire_constant <= "0000000000001000";
    type_cast_1474_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_169_wire_constant <= "0000000000001000";
    type_cast_194_wire_constant <= "0000000000001000";
    type_cast_234_wire_constant <= "00000000000000000000000000000010";
    type_cast_240_wire_constant <= "00000000000000000000000000000001";
    type_cast_246_wire_constant <= "01111111111111111111111111111110";
    type_cast_295_wire_constant <= "0000000000001000";
    type_cast_320_wire_constant <= "0000000000001000";
    type_cast_345_wire_constant <= "0000000000001000";
    type_cast_370_wire_constant <= "0000000000001000";
    type_cast_395_wire_constant <= "0000000000001000";
    type_cast_413_wire_constant <= "00000000000000000000000000000011";
    type_cast_429_wire_constant <= "00000000000000000000000000000011";
    type_cast_442_wire_constant <= "00000000000000000000000000000001";
    type_cast_448_wire_constant <= "11111111111111111111111111111111";
    type_cast_44_wire_constant <= "0000000000001000";
    type_cast_458_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_465_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_474_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_495_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_513_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_531_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_549_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_567_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_585_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_603_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_625_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_643_wire_constant <= "00000000000000000000000000000010";
    type_cast_649_wire_constant <= "00000000000000000000000000000001";
    type_cast_655_wire_constant <= "11111111111111111111111111111111";
    type_cast_665_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_672_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_681_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_69_wire_constant <= "0000000000001000";
    type_cast_702_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_720_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_738_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_756_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_774_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_792_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_810_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_832_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_874_wire_constant <= "00000000000000000000000000000011";
    type_cast_887_wire_constant <= "00000000000000000000000000000010";
    type_cast_893_wire_constant <= "00000000000000000000000000000001";
    type_cast_899_wire_constant <= "11111111111111111111111111111111";
    type_cast_909_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_916_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_927_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_939_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_944_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_94_wire_constant <= "0000000000001000";
    phi_stmt_1354: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1358_wire_constant & type_cast_1360_wire;
      req <= phi_stmt_1354_req_0 & phi_stmt_1354_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1354",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1354_ack_0,
          idata => idata,
          odata => indvar_1354,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1354
    phi_stmt_470: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_474_wire_constant & type_cast_476_wire;
      req <= phi_stmt_470_req_0 & phi_stmt_470_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_470",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_470_ack_0,
          idata => idata,
          odata => indvar556_470,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_470
    phi_stmt_677: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_681_wire_constant & type_cast_683_wire;
      req <= phi_stmt_677_req_0 & phi_stmt_677_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_677",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_677_ack_0,
          idata => idata,
          odata => indvar540_677,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_677
    phi_stmt_921: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_924_wire & type_cast_927_wire_constant;
      req <= phi_stmt_921_req_0 & phi_stmt_921_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_921",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_921_ack_0,
          idata => idata,
          odata => indvar526_921,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_921
    -- flow-through select operator MUX_1350_inst
    tmp525_1351 <= xx_xop_1344 when (tmp522_1328(0) /=  '0') else type_cast_1349_wire_constant;
    -- flow-through select operator MUX_466_inst
    tmp568_467 <= xx_xop572_460 when (tmp564_444(0) /=  '0') else type_cast_465_wire_constant;
    -- flow-through select operator MUX_673_inst
    tmp554_674 <= xx_xop571_667 when (tmp550_651(0) /=  '0') else type_cast_672_wire_constant;
    -- flow-through select operator MUX_917_inst
    tmp538_918 <= xx_xop570_911 when (tmp534_895(0) /=  '0') else type_cast_916_wire_constant;
    addr_of_1367_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1367_final_reg_req_0;
      addr_of_1367_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1367_final_reg_req_1;
      addr_of_1367_final_reg_ack_1<= rack(0);
      addr_of_1367_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1367_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1366_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx433_1368,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_483_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_483_final_reg_req_0;
      addr_of_483_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_483_final_reg_req_1;
      addr_of_483_final_reg_ack_1<= rack(0);
      addr_of_483_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_483_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_482_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_484,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_690_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_690_final_reg_req_0;
      addr_of_690_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_690_final_reg_req_1;
      addr_of_690_final_reg_ack_1<= rack(0);
      addr_of_690_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_690_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 11,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_689_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx246_691,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_934_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_934_final_reg_req_0;
      addr_of_934_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_934_final_reg_req_1;
      addr_of_934_final_reg_ack_1<= rack(0);
      addr_of_934_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_934_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_933_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx269_935,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_102_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_102_inst_req_0;
      type_cast_102_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_102_inst_req_1;
      type_cast_102_inst_ack_1<= rack(0);
      type_cast_102_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_102_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call19_99,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv20_103,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1050_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1050_inst_req_0;
      type_cast_1050_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1050_inst_req_1;
      type_cast_1050_inst_ack_1<= rack(0);
      type_cast_1050_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1050_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr304_1047,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv305_1051,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1057_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1057_inst_req_0;
      type_cast_1057_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1057_inst_req_1;
      type_cast_1057_inst_ack_1<= rack(0);
      type_cast_1057_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1057_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr_236,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv307_1058,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1106_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1106_inst_req_0;
      type_cast_1106_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1106_inst_req_1;
      type_cast_1106_inst_ack_1<= rack(0);
      type_cast_1106_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1106_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr321_1103,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv322_1107,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1113_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1113_inst_req_0;
      type_cast_1113_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1113_inst_req_1;
      type_cast_1113_inst_ack_1<= rack(0);
      type_cast_1113_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1113_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add74_248,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv324_1114,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_114_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_114_inst_req_0;
      type_cast_114_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_114_inst_req_1;
      type_cast_114_inst_ack_1<= rack(0);
      type_cast_114_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_114_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call23_111,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv26_115,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1162_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1162_inst_req_0;
      type_cast_1162_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1162_inst_req_1;
      type_cast_1162_inst_ack_1<= rack(0);
      type_cast_1162_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1162_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr338_1159,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv339_1163,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1169_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1169_inst_req_0;
      type_cast_1169_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1169_inst_req_1;
      type_cast_1169_inst_ack_1<= rack(0);
      type_cast_1169_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1169_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add79_253,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv341_1170,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1201_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1201_inst_req_0;
      type_cast_1201_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1201_inst_req_1;
      type_cast_1201_inst_ack_1<= rack(0);
      type_cast_1201_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1201_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1200_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv355_1202,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1213_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1213_inst_req_0;
      type_cast_1213_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1213_inst_req_1;
      type_cast_1213_inst_ack_1<= rack(0);
      type_cast_1213_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1213_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub_1207,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv362_1214,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1223_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1223_inst_req_0;
      type_cast_1223_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1223_inst_req_1;
      type_cast_1223_inst_ack_1<= rack(0);
      type_cast_1223_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1223_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr365_1220,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv368_1224,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1233_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1233_inst_req_0;
      type_cast_1233_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1233_inst_req_1;
      type_cast_1233_inst_ack_1<= rack(0);
      type_cast_1233_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1233_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr371_1230,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv374_1234,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1243_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1243_inst_req_0;
      type_cast_1243_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1243_inst_req_1;
      type_cast_1243_inst_ack_1<= rack(0);
      type_cast_1243_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1243_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr377_1240,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv380_1244,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1253_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1253_inst_req_0;
      type_cast_1253_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1253_inst_req_1;
      type_cast_1253_inst_ack_1<= rack(0);
      type_cast_1253_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1253_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr383_1250,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv386_1254,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1263_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1263_inst_req_0;
      type_cast_1263_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1263_inst_req_1;
      type_cast_1263_inst_ack_1<= rack(0);
      type_cast_1263_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1263_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr389_1260,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv392_1264,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1273_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1273_inst_req_0;
      type_cast_1273_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1273_inst_req_1;
      type_cast_1273_inst_ack_1<= rack(0);
      type_cast_1273_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1273_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr395_1270,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv398_1274,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_127_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_127_inst_req_0;
      type_cast_127_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_127_inst_req_1;
      type_cast_127_inst_ack_1<= rack(0);
      type_cast_127_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_127_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call28_124,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_128,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1283_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1283_inst_req_0;
      type_cast_1283_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1283_inst_req_1;
      type_cast_1283_inst_ack_1<= rack(0);
      type_cast_1283_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1283_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr401_1280,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv404_1284,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1337_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1337_inst_req_0;
      type_cast_1337_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1337_inst_req_1;
      type_cast_1337_inst_ack_1<= rack(0);
      type_cast_1337_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1337_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp521x_xop_1334,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_197_1338,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1360_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1360_inst_req_0;
      type_cast_1360_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1360_inst_req_1;
      type_cast_1360_inst_ack_1<= rack(0);
      type_cast_1360_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1360_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1476,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1360_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1375_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1375_inst_req_0;
      type_cast_1375_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1375_inst_req_1;
      type_cast_1375_inst_ack_1<= rack(0);
      type_cast_1375_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1375_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp434_1372,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv438_1376,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1385_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1385_inst_req_0;
      type_cast_1385_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1385_inst_req_1;
      type_cast_1385_inst_ack_1<= rack(0);
      type_cast_1385_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1385_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr441_1382,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv444_1386,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1395_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1395_inst_req_0;
      type_cast_1395_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1395_inst_req_1;
      type_cast_1395_inst_ack_1<= rack(0);
      type_cast_1395_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1395_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr447_1392,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv450_1396,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_139_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_139_inst_req_0;
      type_cast_139_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_139_inst_req_1;
      type_cast_139_inst_ack_1<= rack(0);
      type_cast_139_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_139_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call32_136,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv35_140,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1405_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1405_inst_req_0;
      type_cast_1405_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1405_inst_req_1;
      type_cast_1405_inst_ack_1<= rack(0);
      type_cast_1405_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1405_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr453_1402,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv456_1406,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1415_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1415_inst_req_0;
      type_cast_1415_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1415_inst_req_1;
      type_cast_1415_inst_ack_1<= rack(0);
      type_cast_1415_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1415_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr459_1412,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv462_1416,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1425_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1425_inst_req_0;
      type_cast_1425_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1425_inst_req_1;
      type_cast_1425_inst_ack_1<= rack(0);
      type_cast_1425_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1425_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr465_1422,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv468_1426,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1435_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1435_inst_req_0;
      type_cast_1435_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1435_inst_req_1;
      type_cast_1435_inst_ack_1<= rack(0);
      type_cast_1435_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1435_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr471_1432,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv474_1436,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1445_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1445_inst_req_0;
      type_cast_1445_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1445_inst_req_1;
      type_cast_1445_inst_ack_1<= rack(0);
      type_cast_1445_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1445_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr477_1442,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv480_1446,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_152_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_152_inst_req_0;
      type_cast_152_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_152_inst_req_1;
      type_cast_152_inst_ack_1<= rack(0);
      type_cast_152_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_152_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call37_149,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_153,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_164_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_164_inst_req_0;
      type_cast_164_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_164_inst_req_1;
      type_cast_164_inst_ack_1<= rack(0);
      type_cast_164_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_164_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_161,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_165,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_177_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_177_inst_req_0;
      type_cast_177_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_177_inst_req_1;
      type_cast_177_inst_ack_1<= rack(0);
      type_cast_177_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_177_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_174,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv47_178,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_189_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_189_inst_req_0;
      type_cast_189_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_189_inst_req_1;
      type_cast_189_inst_ack_1<= rack(0);
      type_cast_189_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_189_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call50_186,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv53_190,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_202_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_202_inst_req_0;
      type_cast_202_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_202_inst_req_1;
      type_cast_202_inst_ack_1<= rack(0);
      type_cast_202_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_202_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call55_199,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_203,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_211_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_211_inst_req_0;
      type_cast_211_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_211_inst_req_1;
      type_cast_211_inst_ack_1<= rack(0);
      type_cast_211_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_211_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_58,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv61_212,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_215_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_215_inst_req_0;
      type_cast_215_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_215_inst_req_1;
      type_cast_215_inst_ack_1<= rack(0);
      type_cast_215_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_215_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add12_83,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv63_216,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_219_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_219_inst_req_0;
      type_cast_219_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_219_inst_req_1;
      type_cast_219_inst_ack_1<= rack(0);
      type_cast_219_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_219_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add21_108,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_220,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_256_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_256_inst_req_0;
      type_cast_256_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_256_inst_req_1;
      type_cast_256_inst_ack_1<= rack(0);
      type_cast_256_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_256_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add30_133,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv82_257,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_260_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_260_inst_req_0;
      type_cast_260_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_260_inst_req_1;
      type_cast_260_inst_ack_1<= rack(0);
      type_cast_260_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_260_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add39_158,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv84_261,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_264_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_264_inst_req_0;
      type_cast_264_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_264_inst_req_1;
      type_cast_264_inst_ack_1<= rack(0);
      type_cast_264_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_264_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add48_183,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv87_265,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_268_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_268_inst_req_0;
      type_cast_268_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_268_inst_req_1;
      type_cast_268_inst_ack_1<= rack(0);
      type_cast_268_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_268_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add57_208,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_269,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_290_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_290_inst_req_0;
      type_cast_290_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_290_inst_req_1;
      type_cast_290_inst_ack_1<= rack(0);
      type_cast_290_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_290_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call92_287,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_291,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_303_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_303_inst_req_0;
      type_cast_303_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_303_inst_req_1;
      type_cast_303_inst_ack_1<= rack(0);
      type_cast_303_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_303_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call97_300,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv98_304,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_315_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_315_inst_req_0;
      type_cast_315_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_315_inst_req_1;
      type_cast_315_inst_ack_1<= rack(0);
      type_cast_315_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_315_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call101_312,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv104_316,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_328_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_328_inst_req_0;
      type_cast_328_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_328_inst_req_1;
      type_cast_328_inst_ack_1<= rack(0);
      type_cast_328_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_328_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call106_325,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv107_329,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_340_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_340_inst_req_0;
      type_cast_340_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_340_inst_req_1;
      type_cast_340_inst_ack_1<= rack(0);
      type_cast_340_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_340_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call110_337,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv113_341,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_353_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_353_inst_req_0;
      type_cast_353_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_353_inst_req_1;
      type_cast_353_inst_ack_1<= rack(0);
      type_cast_353_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_353_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call115_350,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv116_354,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_365_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_365_inst_req_0;
      type_cast_365_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_365_inst_req_1;
      type_cast_365_inst_ack_1<= rack(0);
      type_cast_365_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_365_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call119_362,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv122_366,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_378_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_378_inst_req_0;
      type_cast_378_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_378_inst_req_1;
      type_cast_378_inst_ack_1<= rack(0);
      type_cast_378_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_378_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call124_375,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv125_379,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_390_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_390_inst_req_0;
      type_cast_390_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_390_inst_req_1;
      type_cast_390_inst_ack_1<= rack(0);
      type_cast_390_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_390_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call128_387,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv131_391,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_39_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_39_inst_req_0;
      type_cast_39_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_39_inst_req_1;
      type_cast_39_inst_ack_1<= rack(0);
      type_cast_39_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_39_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_36,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1_40,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_403_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_403_inst_req_0;
      type_cast_403_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_403_inst_req_1;
      type_cast_403_inst_ack_1<= rack(0);
      type_cast_403_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_403_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call133_400,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv134_404,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_453_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_453_inst_req_0;
      type_cast_453_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_453_inst_req_1;
      type_cast_453_inst_ack_1<= rack(0);
      type_cast_453_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_453_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp563x_xop_450,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_26_454,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_476_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_476_inst_req_0;
      type_cast_476_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_476_inst_req_1;
      type_cast_476_inst_ack_1<= rack(0);
      type_cast_476_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_476_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext557_627,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_476_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_490_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_490_inst_req_0;
      type_cast_490_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_490_inst_req_1;
      type_cast_490_inst_ack_1<= rack(0);
      type_cast_490_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_490_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call143_487,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv144_491,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_503_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_503_inst_req_0;
      type_cast_503_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_503_inst_req_1;
      type_cast_503_inst_ack_1<= rack(0);
      type_cast_503_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_503_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call147_500,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv149_504,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_521_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_521_inst_req_0;
      type_cast_521_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_521_inst_req_1;
      type_cast_521_inst_ack_1<= rack(0);
      type_cast_521_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_521_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call153_518,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv155_522,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_52_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_52_inst_req_0;
      type_cast_52_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_52_inst_req_1;
      type_cast_52_inst_ack_1<= rack(0);
      type_cast_52_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_52_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_49,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_53,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_539_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_539_inst_req_0;
      type_cast_539_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_539_inst_req_1;
      type_cast_539_inst_ack_1<= rack(0);
      type_cast_539_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_539_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call159_536,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv161_540,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_557_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_557_inst_req_0;
      type_cast_557_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_557_inst_req_1;
      type_cast_557_inst_ack_1<= rack(0);
      type_cast_557_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_557_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call165_554,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv167_558,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_575_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_575_inst_req_0;
      type_cast_575_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_575_inst_req_1;
      type_cast_575_inst_ack_1<= rack(0);
      type_cast_575_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_575_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call171_572,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv173_576,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_593_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_593_inst_req_0;
      type_cast_593_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_593_inst_req_1;
      type_cast_593_inst_ack_1<= rack(0);
      type_cast_593_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_593_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call177_590,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv179_594,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_611_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_611_inst_req_0;
      type_cast_611_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_611_inst_req_1;
      type_cast_611_inst_ack_1<= rack(0);
      type_cast_611_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_611_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call183_608,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv185_612,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_64_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_64_inst_req_0;
      type_cast_64_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_64_inst_req_1;
      type_cast_64_inst_ack_1<= rack(0);
      type_cast_64_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_64_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_61,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv8_65,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_660_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_660_inst_req_0;
      type_cast_660_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_660_inst_req_1;
      type_cast_660_inst_ack_1<= rack(0);
      type_cast_660_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_660_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp549x_xop_657,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_39_661,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_683_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_683_inst_req_0;
      type_cast_683_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_683_inst_req_1;
      type_cast_683_inst_ack_1<= rack(0);
      type_cast_683_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_683_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext541_834,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_683_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_697_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_697_inst_req_0;
      type_cast_697_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_697_inst_req_1;
      type_cast_697_inst_ack_1<= rack(0);
      type_cast_697_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_697_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call199_694,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv200_698,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_710_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_710_inst_req_0;
      type_cast_710_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_710_inst_req_1;
      type_cast_710_inst_ack_1<= rack(0);
      type_cast_710_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_710_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call203_707,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv205_711,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_728_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_728_inst_req_0;
      type_cast_728_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_728_inst_req_1;
      type_cast_728_inst_ack_1<= rack(0);
      type_cast_728_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_728_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call209_725,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv211_729,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_746_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_746_inst_req_0;
      type_cast_746_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_746_inst_req_1;
      type_cast_746_inst_ack_1<= rack(0);
      type_cast_746_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_746_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call215_743,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv217_747,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_764_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_764_inst_req_0;
      type_cast_764_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_764_inst_req_1;
      type_cast_764_inst_ack_1<= rack(0);
      type_cast_764_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_764_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call221_761,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv223_765,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_77_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_77_inst_req_0;
      type_cast_77_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_77_inst_req_1;
      type_cast_77_inst_ack_1<= rack(0);
      type_cast_77_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_77_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call10_74,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv11_78,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_782_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_782_inst_req_0;
      type_cast_782_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_782_inst_req_1;
      type_cast_782_inst_ack_1<= rack(0);
      type_cast_782_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_782_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call227_779,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv229_783,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_800_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_800_inst_req_0;
      type_cast_800_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_800_inst_req_1;
      type_cast_800_inst_ack_1<= rack(0);
      type_cast_800_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_800_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call233_797,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv235_801,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_818_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_818_inst_req_0;
      type_cast_818_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_818_inst_req_1;
      type_cast_818_inst_ack_1<= rack(0);
      type_cast_818_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_818_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call239_815,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv241_819,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_851_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_851_inst_req_0;
      type_cast_851_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_851_inst_req_1;
      type_cast_851_inst_ack_1<= rack(0);
      type_cast_851_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_851_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add117_359,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv253_852,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_855_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_855_inst_req_0;
      type_cast_855_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_855_inst_req_1;
      type_cast_855_inst_ack_1<= rack(0);
      type_cast_855_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_855_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add126_384,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv255_856,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_859_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_859_inst_req_0;
      type_cast_859_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_859_inst_req_1;
      type_cast_859_inst_ack_1<= rack(0);
      type_cast_859_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_859_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add135_409,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv258_860,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_89_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_89_inst_req_0;
      type_cast_89_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_89_inst_req_1;
      type_cast_89_inst_ack_1<= rack(0);
      type_cast_89_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_89_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call14_86,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_90,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_904_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_904_inst_req_0;
      type_cast_904_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_904_inst_req_1;
      type_cast_904_inst_ack_1<= rack(0);
      type_cast_904_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_904_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp533x_xop_901,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_53_905,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_924_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_924_inst_req_0;
      type_cast_924_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_924_inst_req_1;
      type_cast_924_inst_ack_1<= rack(0);
      type_cast_924_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_924_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext527_946,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_924_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_968_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_968_inst_req_0;
      type_cast_968_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_968_inst_req_1;
      type_cast_968_inst_ack_1<= rack(0);
      type_cast_968_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_968_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_967_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv276_969,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1366_index_1_rename
    process(R_indvar_1365_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_1365_resized;
      ov(13 downto 0) := iv;
      R_indvar_1365_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1366_index_1_resize
    process(indvar_1354) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_1354;
      ov := iv(13 downto 0);
      R_indvar_1365_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1366_root_address_inst
    process(array_obj_ref_1366_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1366_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1366_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_482_index_1_rename
    process(R_indvar556_481_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar556_481_resized;
      ov(13 downto 0) := iv;
      R_indvar556_481_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_482_index_1_resize
    process(indvar556_470) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar556_470;
      ov := iv(13 downto 0);
      R_indvar556_481_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_482_root_address_inst
    process(array_obj_ref_482_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_482_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_482_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_689_index_1_rename
    process(R_indvar540_688_resized) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar540_688_resized;
      ov(10 downto 0) := iv;
      R_indvar540_688_scaled <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_689_index_1_resize
    process(indvar540_677) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar540_677;
      ov := iv(10 downto 0);
      R_indvar540_688_resized <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_689_root_address_inst
    process(array_obj_ref_689_final_offset) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_689_final_offset;
      ov(10 downto 0) := iv;
      array_obj_ref_689_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_933_index_1_rename
    process(R_indvar526_932_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar526_932_resized;
      ov(13 downto 0) := iv;
      R_indvar526_932_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_933_index_1_resize
    process(indvar526_921) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar526_921;
      ov := iv(13 downto 0);
      R_indvar526_932_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_933_root_address_inst
    process(array_obj_ref_933_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_933_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_933_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1371_addr_0
    process(ptr_deref_1371_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1371_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1371_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1371_base_resize
    process(arrayidx433_1368) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx433_1368;
      ov := iv(13 downto 0);
      ptr_deref_1371_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1371_gather_scatter
    process(ptr_deref_1371_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1371_data_0;
      ov(63 downto 0) := iv;
      tmp434_1372 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1371_root_address_inst
    process(ptr_deref_1371_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1371_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1371_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_619_addr_0
    process(ptr_deref_619_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_619_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_619_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_619_base_resize
    process(arrayidx_484) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_484;
      ov := iv(13 downto 0);
      ptr_deref_619_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_619_gather_scatter
    process(add186_617) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add186_617;
      ov(63 downto 0) := iv;
      ptr_deref_619_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_619_root_address_inst
    process(ptr_deref_619_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_619_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_619_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_826_addr_0
    process(ptr_deref_826_root_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_826_root_address;
      ov(10 downto 0) := iv;
      ptr_deref_826_word_address_0 <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_826_base_resize
    process(arrayidx246_691) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx246_691;
      ov := iv(10 downto 0);
      ptr_deref_826_resized_base_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_826_gather_scatter
    process(add242_824) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add242_824;
      ov(63 downto 0) := iv;
      ptr_deref_826_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_826_root_address_inst
    process(ptr_deref_826_resized_base_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_826_resized_base_address;
      ov(10 downto 0) := iv;
      ptr_deref_826_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_937_addr_0
    process(ptr_deref_937_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_937_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_937_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_937_base_resize
    process(arrayidx269_935) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx269_935;
      ov := iv(13 downto 0);
      ptr_deref_937_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_937_gather_scatter
    process(type_cast_939_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_939_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_937_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_937_root_address_inst
    process(ptr_deref_937_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_937_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_937_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1310_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp264506_876;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1310_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1310_branch_req_0,
          ack0 => if_stmt_1310_branch_ack_0,
          ack1 => if_stmt_1310_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1482_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_1481;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1482_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1482_branch_req_0,
          ack0 => if_stmt_1482_branch_ack_0,
          ack1 => if_stmt_1482_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_417_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp514_416;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_417_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_417_branch_req_0,
          ack0 => if_stmt_417_branch_ack_0,
          ack1 => if_stmt_417_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_432_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp194510_431;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_432_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_432_branch_req_0,
          ack0 => if_stmt_432_branch_ack_0,
          ack1 => if_stmt_432_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_633_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond3_632;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_633_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_633_branch_req_0,
          ack0 => if_stmt_633_branch_ack_0,
          ack1 => if_stmt_633_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_840_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond2_839;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_840_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_840_branch_req_0,
          ack0 => if_stmt_840_branch_ack_0,
          ack1 => if_stmt_840_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_877_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp264506_876;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_877_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_877_branch_req_0,
          ack0 => if_stmt_877_branch_ack_0,
          ack1 => if_stmt_877_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_952_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_951;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_952_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_952_branch_req_0,
          ack0 => if_stmt_952_branch_ack_0,
          ack1 => if_stmt_952_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_1333_inst
    process(tmp521_1322) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp521_1322, type_cast_1332_wire_constant, tmp_var);
      tmp521x_xop_1334 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_252_inst
    process(add74_248, shr_236) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add74_248, shr_236, tmp_var);
      add79_253 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_449_inst
    process(shr_236) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr_236, type_cast_448_wire_constant, tmp_var);
      tmp563x_xop_450 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_656_inst
    process(tmp549_645) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp549_645, type_cast_655_wire_constant, tmp_var);
      tmp549x_xop_657 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_900_inst
    process(tmp533_889) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp533_889, type_cast_899_wire_constant, tmp_var);
      tmp533x_xop_901 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1343_inst
    process(iNsTr_197_1338) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_197_1338, type_cast_1342_wire_constant, tmp_var);
      xx_xop_1344 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1475_inst
    process(indvar_1354) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1354, type_cast_1474_wire_constant, tmp_var);
      indvarx_xnext_1476 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_459_inst
    process(iNsTr_26_454) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_26_454, type_cast_458_wire_constant, tmp_var);
      xx_xop572_460 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_626_inst
    process(indvar556_470) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar556_470, type_cast_625_wire_constant, tmp_var);
      indvarx_xnext557_627 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_666_inst
    process(iNsTr_39_661) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_39_661, type_cast_665_wire_constant, tmp_var);
      xx_xop571_667 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_833_inst
    process(indvar540_677) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar540_677, type_cast_832_wire_constant, tmp_var);
      indvarx_xnext541_834 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_910_inst
    process(iNsTr_53_905) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_53_905, type_cast_909_wire_constant, tmp_var);
      xx_xop570_911 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_945_inst
    process(indvar526_921) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar526_921, type_cast_944_wire_constant, tmp_var);
      indvarx_xnext527_946 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_247_inst
    process(iNsTr_14_242) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(iNsTr_14_242, type_cast_246_wire_constant, tmp_var);
      add74_248 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1480_inst
    process(indvarx_xnext_1476, tmp525_1351) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1476, tmp525_1351, tmp_var);
      exitcond1_1481 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_631_inst
    process(indvarx_xnext557_627, tmp568_467) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext557_627, tmp568_467, tmp_var);
      exitcond3_632 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_838_inst
    process(indvarx_xnext541_834, tmp554_674) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext541_834, tmp554_674, tmp_var);
      exitcond2_839 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_950_inst
    process(indvarx_xnext527_946, tmp538_918) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext527_946, tmp538_918, tmp_var);
      exitcond_951 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1046_inst
    process(mul66_230) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_230, type_cast_1045_wire_constant, tmp_var);
      shr304_1047 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1102_inst
    process(mul66_230) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_230, type_cast_1101_wire_constant, tmp_var);
      shr321_1103 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1158_inst
    process(add79_253) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add79_253, type_cast_1157_wire_constant, tmp_var);
      shr338_1159 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1321_inst
    process(mul259_870) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul259_870, type_cast_1320_wire_constant, tmp_var);
      tmp521_1322 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_235_inst
    process(mul66_230) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_230, type_cast_234_wire_constant, tmp_var);
      shr_236 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_241_inst
    process(mul66_230) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_230, type_cast_240_wire_constant, tmp_var);
      iNsTr_14_242 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_644_inst
    process(mul91_284) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul91_284, type_cast_643_wire_constant, tmp_var);
      tmp549_645 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_888_inst
    process(mul259_870) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul259_870, type_cast_887_wire_constant, tmp_var);
      tmp533_889 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1219_inst
    process(sub_1207) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1207, type_cast_1218_wire_constant, tmp_var);
      shr365_1220 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1229_inst
    process(sub_1207) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1207, type_cast_1228_wire_constant, tmp_var);
      shr371_1230 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1239_inst
    process(sub_1207) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1207, type_cast_1238_wire_constant, tmp_var);
      shr377_1240 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1249_inst
    process(sub_1207) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1207, type_cast_1248_wire_constant, tmp_var);
      shr383_1250 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1259_inst
    process(sub_1207) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1207, type_cast_1258_wire_constant, tmp_var);
      shr389_1260 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1269_inst
    process(sub_1207) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1207, type_cast_1268_wire_constant, tmp_var);
      shr395_1270 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1279_inst
    process(sub_1207) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1207, type_cast_1278_wire_constant, tmp_var);
      shr401_1280 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1381_inst
    process(tmp434_1372) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp434_1372, type_cast_1380_wire_constant, tmp_var);
      shr441_1382 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1391_inst
    process(tmp434_1372) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp434_1372, type_cast_1390_wire_constant, tmp_var);
      shr447_1392 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1401_inst
    process(tmp434_1372) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp434_1372, type_cast_1400_wire_constant, tmp_var);
      shr453_1402 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1411_inst
    process(tmp434_1372) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp434_1372, type_cast_1410_wire_constant, tmp_var);
      shr459_1412 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1421_inst
    process(tmp434_1372) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp434_1372, type_cast_1420_wire_constant, tmp_var);
      shr465_1422 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1431_inst
    process(tmp434_1372) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp434_1372, type_cast_1430_wire_constant, tmp_var);
      shr471_1432 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1441_inst
    process(tmp434_1372) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp434_1372, type_cast_1440_wire_constant, tmp_var);
      shr477_1442 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_224_inst
    process(conv63_216, conv61_212) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv63_216, conv61_212, tmp_var);
      mul_225 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_229_inst
    process(mul_225, conv65_220) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_225, conv65_220, tmp_var);
      mul66_230 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_273_inst
    process(conv84_261, conv82_257) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv84_261, conv82_257, tmp_var);
      mul85_274 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_278_inst
    process(mul85_274, conv87_265) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul85_274, conv87_265, tmp_var);
      mul88_279 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_283_inst
    process(mul88_279, conv90_269) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul88_279, conv90_269, tmp_var);
      mul91_284 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_864_inst
    process(conv255_856, conv253_852) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv255_856, conv253_852, tmp_var);
      mul256_865 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_869_inst
    process(mul256_865, conv258_860) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul256_865, conv258_860, tmp_var);
      mul259_870 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_107_inst
    process(shl18_96, conv20_103) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl18_96, conv20_103, tmp_var);
      add21_108 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_132_inst
    process(shl27_121, conv29_128) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl27_121, conv29_128, tmp_var);
      add30_133 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_157_inst
    process(shl36_146, conv38_153) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl36_146, conv38_153, tmp_var);
      add39_158 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_182_inst
    process(shl45_171, conv47_178) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl45_171, conv47_178, tmp_var);
      add48_183 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_207_inst
    process(shl54_196, conv56_203) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl54_196, conv56_203, tmp_var);
      add57_208 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_308_inst
    process(shl96_297, conv98_304) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl96_297, conv98_304, tmp_var);
      add99_309 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_333_inst
    process(shl105_322, conv107_329) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl105_322, conv107_329, tmp_var);
      add108_334 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_358_inst
    process(shl114_347, conv116_354) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl114_347, conv116_354, tmp_var);
      add117_359 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_383_inst
    process(shl123_372, conv125_379) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl123_372, conv125_379, tmp_var);
      add126_384 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_408_inst
    process(shl132_397, conv134_404) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl132_397, conv134_404, tmp_var);
      add135_409 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_57_inst
    process(shl_46, conv3_53) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_46, conv3_53, tmp_var);
      add_58 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_82_inst
    process(shl9_71, conv11_78) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl9_71, conv11_78, tmp_var);
      add12_83 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_508_inst
    process(shl146_497, conv149_504) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl146_497, conv149_504, tmp_var);
      add150_509 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_526_inst
    process(shl152_515, conv155_522) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl152_515, conv155_522, tmp_var);
      add156_527 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_544_inst
    process(shl158_533, conv161_540) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl158_533, conv161_540, tmp_var);
      add162_545 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_562_inst
    process(shl164_551, conv167_558) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl164_551, conv167_558, tmp_var);
      add168_563 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_580_inst
    process(shl170_569, conv173_576) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl170_569, conv173_576, tmp_var);
      add174_581 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_598_inst
    process(shl176_587, conv179_594) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl176_587, conv179_594, tmp_var);
      add180_599 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_616_inst
    process(shl182_605, conv185_612) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl182_605, conv185_612, tmp_var);
      add186_617 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_715_inst
    process(shl202_704, conv205_711) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl202_704, conv205_711, tmp_var);
      add206_716 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_733_inst
    process(shl208_722, conv211_729) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl208_722, conv211_729, tmp_var);
      add212_734 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_751_inst
    process(shl214_740, conv217_747) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl214_740, conv217_747, tmp_var);
      add218_752 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_769_inst
    process(shl220_758, conv223_765) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl220_758, conv223_765, tmp_var);
      add224_770 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_787_inst
    process(shl226_776, conv229_783) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl226_776, conv229_783, tmp_var);
      add230_788 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_805_inst
    process(shl232_794, conv235_801) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl232_794, conv235_801, tmp_var);
      add236_806 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_823_inst
    process(shl238_812, conv241_819) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl238_812, conv241_819, tmp_var);
      add242_824 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_120_inst
    process(conv26_115) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv26_115, type_cast_119_wire_constant, tmp_var);
      shl27_121 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_145_inst
    process(conv35_140) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv35_140, type_cast_144_wire_constant, tmp_var);
      shl36_146 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_170_inst
    process(conv44_165) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv44_165, type_cast_169_wire_constant, tmp_var);
      shl45_171 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_195_inst
    process(conv53_190) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv53_190, type_cast_194_wire_constant, tmp_var);
      shl54_196 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_296_inst
    process(conv95_291) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv95_291, type_cast_295_wire_constant, tmp_var);
      shl96_297 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_321_inst
    process(conv104_316) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv104_316, type_cast_320_wire_constant, tmp_var);
      shl105_322 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_346_inst
    process(conv113_341) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv113_341, type_cast_345_wire_constant, tmp_var);
      shl114_347 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_371_inst
    process(conv122_366) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv122_366, type_cast_370_wire_constant, tmp_var);
      shl123_372 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_396_inst
    process(conv131_391) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv131_391, type_cast_395_wire_constant, tmp_var);
      shl132_397 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_45_inst
    process(conv1_40) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1_40, type_cast_44_wire_constant, tmp_var);
      shl_46 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_70_inst
    process(conv8_65) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv8_65, type_cast_69_wire_constant, tmp_var);
      shl9_71 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_95_inst
    process(conv17_90) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv17_90, type_cast_94_wire_constant, tmp_var);
      shl18_96 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_496_inst
    process(conv144_491) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv144_491, type_cast_495_wire_constant, tmp_var);
      shl146_497 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_514_inst
    process(add150_509) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add150_509, type_cast_513_wire_constant, tmp_var);
      shl152_515 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_532_inst
    process(add156_527) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add156_527, type_cast_531_wire_constant, tmp_var);
      shl158_533 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_550_inst
    process(add162_545) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add162_545, type_cast_549_wire_constant, tmp_var);
      shl164_551 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_568_inst
    process(add168_563) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add168_563, type_cast_567_wire_constant, tmp_var);
      shl170_569 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_586_inst
    process(add174_581) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add174_581, type_cast_585_wire_constant, tmp_var);
      shl176_587 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_604_inst
    process(add180_599) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add180_599, type_cast_603_wire_constant, tmp_var);
      shl182_605 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_703_inst
    process(conv200_698) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv200_698, type_cast_702_wire_constant, tmp_var);
      shl202_704 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_721_inst
    process(add206_716) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add206_716, type_cast_720_wire_constant, tmp_var);
      shl208_722 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_739_inst
    process(add212_734) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add212_734, type_cast_738_wire_constant, tmp_var);
      shl214_740 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_757_inst
    process(add218_752) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add218_752, type_cast_756_wire_constant, tmp_var);
      shl220_758 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_775_inst
    process(add224_770) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add224_770, type_cast_774_wire_constant, tmp_var);
      shl226_776 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_793_inst
    process(add230_788) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add230_788, type_cast_792_wire_constant, tmp_var);
      shl232_794 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_811_inst
    process(add236_806) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add236_806, type_cast_810_wire_constant, tmp_var);
      shl238_812 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_1206_inst
    process(conv355_1202, conv276_969) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv355_1202, conv276_969, tmp_var);
      sub_1207 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1327_inst
    process(tmp521_1322) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp521_1322, type_cast_1326_wire_constant, tmp_var);
      tmp522_1328 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_414_inst
    process(mul66_230) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul66_230, type_cast_413_wire_constant, tmp_var);
      cmp514_416 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_430_inst
    process(mul91_284) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul91_284, type_cast_429_wire_constant, tmp_var);
      cmp194510_431 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_443_inst
    process(shr_236) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(shr_236, type_cast_442_wire_constant, tmp_var);
      tmp564_444 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_650_inst
    process(tmp549_645) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp549_645, type_cast_649_wire_constant, tmp_var);
      tmp550_651 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_875_inst
    process(mul259_870) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul259_870, type_cast_874_wire_constant, tmp_var);
      cmp264506_876 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_894_inst
    process(tmp533_889) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp533_889, type_cast_893_wire_constant, tmp_var);
      tmp534_895 <= tmp_var; --
    end process;
    -- shared split operator group (107) : array_obj_ref_1366_index_offset 
    ApIntAdd_group_107: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_1365_scaled;
      array_obj_ref_1366_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1366_index_offset_req_0;
      array_obj_ref_1366_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1366_index_offset_req_1;
      array_obj_ref_1366_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_107_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_107_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_107",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 107
    -- shared split operator group (108) : array_obj_ref_482_index_offset 
    ApIntAdd_group_108: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar556_481_scaled;
      array_obj_ref_482_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_482_index_offset_req_0;
      array_obj_ref_482_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_482_index_offset_req_1;
      array_obj_ref_482_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_108_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_108_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_108",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 108
    -- shared split operator group (109) : array_obj_ref_689_index_offset 
    ApIntAdd_group_109: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar540_688_scaled;
      array_obj_ref_689_final_offset <= data_out(10 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_689_index_offset_req_0;
      array_obj_ref_689_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_689_index_offset_req_1;
      array_obj_ref_689_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_109_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_109_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_109",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000100010",
          constant_width => 11,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 109
    -- shared split operator group (110) : array_obj_ref_933_index_offset 
    ApIntAdd_group_110: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar526_932_scaled;
      array_obj_ref_933_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_933_index_offset_req_0;
      array_obj_ref_933_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_933_index_offset_req_1;
      array_obj_ref_933_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_110_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_110_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_110",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 110
    -- unary operator type_cast_1200_inst
    process(call354_1197) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call354_1197, tmp_var);
      type_cast_1200_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_967_inst
    process(call275_963) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call275_963, tmp_var);
      type_cast_967_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_1371_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1371_load_0_req_0;
      ptr_deref_1371_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1371_load_0_req_1;
      ptr_deref_1371_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1371_word_address_0;
      ptr_deref_1371_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(13 downto 0),
          mtag => memory_space_3_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(63 downto 0),
          mtag => memory_space_3_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_619_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_619_store_0_req_0;
      ptr_deref_619_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_619_store_0_req_1;
      ptr_deref_619_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_619_word_address_0;
      data_in <= ptr_deref_619_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_826_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(10 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_826_store_0_req_0;
      ptr_deref_826_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_826_store_0_req_1;
      ptr_deref_826_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_826_word_address_0;
      data_in <= ptr_deref_826_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 11,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(10 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_937_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_937_store_0_req_0;
      ptr_deref_937_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_937_store_0_req_1;
      ptr_deref_937_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_937_word_address_0;
      data_in <= ptr_deref_937_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared inport operator group (0) : RPIPE_Block0_done_1184_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block0_done_1184_inst_req_0;
      RPIPE_Block0_done_1184_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block0_done_1184_inst_req_1;
      RPIPE_Block0_done_1184_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call346_1185 <= data_out(15 downto 0);
      Block0_done_read_0_gI: SplitGuardInterface generic map(name => "Block0_done_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_done_read_0: InputPortRevised -- 
        generic map ( name => "Block0_done_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_done_pipe_read_req(0),
          oack => Block0_done_pipe_read_ack(0),
          odata => Block0_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_Block1_done_1187_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block1_done_1187_inst_req_0;
      RPIPE_Block1_done_1187_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block1_done_1187_inst_req_1;
      RPIPE_Block1_done_1187_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call348_1188 <= data_out(15 downto 0);
      Block1_done_read_1_gI: SplitGuardInterface generic map(name => "Block1_done_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_done_read_1: InputPortRevised -- 
        generic map ( name => "Block1_done_read_1", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_done_pipe_read_req(0),
          oack => Block1_done_pipe_read_ack(0),
          odata => Block1_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_Block2_done_1190_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block2_done_1190_inst_req_0;
      RPIPE_Block2_done_1190_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block2_done_1190_inst_req_1;
      RPIPE_Block2_done_1190_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call350_1191 <= data_out(15 downto 0);
      Block2_done_read_2_gI: SplitGuardInterface generic map(name => "Block2_done_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_done_read_2: InputPortRevised -- 
        generic map ( name => "Block2_done_read_2", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_done_pipe_read_req(0),
          oack => Block2_done_pipe_read_ack(0),
          odata => Block2_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_Block3_done_1193_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block3_done_1193_inst_req_0;
      RPIPE_Block3_done_1193_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block3_done_1193_inst_req_1;
      RPIPE_Block3_done_1193_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call352_1194 <= data_out(15 downto 0);
      Block3_done_read_3_gI: SplitGuardInterface generic map(name => "Block3_done_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_done_read_3: InputPortRevised -- 
        generic map ( name => "Block3_done_read_3", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_done_pipe_read_req(0),
          oack => Block3_done_pipe_read_ack(0),
          odata => Block3_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared inport operator group (4) : RPIPE_ConvTranspose_input_pipe_724_inst RPIPE_ConvTranspose_input_pipe_589_inst RPIPE_ConvTranspose_input_pipe_517_inst RPIPE_ConvTranspose_input_pipe_607_inst RPIPE_ConvTranspose_input_pipe_110_inst RPIPE_ConvTranspose_input_pipe_73_inst RPIPE_ConvTranspose_input_pipe_135_inst RPIPE_ConvTranspose_input_pipe_98_inst RPIPE_ConvTranspose_input_pipe_486_inst RPIPE_ConvTranspose_input_pipe_571_inst RPIPE_ConvTranspose_input_pipe_742_inst RPIPE_ConvTranspose_input_pipe_123_inst RPIPE_ConvTranspose_input_pipe_48_inst RPIPE_ConvTranspose_input_pipe_814_inst RPIPE_ConvTranspose_input_pipe_693_inst RPIPE_ConvTranspose_input_pipe_60_inst RPIPE_ConvTranspose_input_pipe_85_inst RPIPE_ConvTranspose_input_pipe_760_inst RPIPE_ConvTranspose_input_pipe_535_inst RPIPE_ConvTranspose_input_pipe_778_inst RPIPE_ConvTranspose_input_pipe_35_inst RPIPE_ConvTranspose_input_pipe_499_inst RPIPE_ConvTranspose_input_pipe_553_inst RPIPE_ConvTranspose_input_pipe_706_inst RPIPE_ConvTranspose_input_pipe_796_inst RPIPE_ConvTranspose_input_pipe_148_inst RPIPE_ConvTranspose_input_pipe_160_inst RPIPE_ConvTranspose_input_pipe_173_inst RPIPE_ConvTranspose_input_pipe_185_inst RPIPE_ConvTranspose_input_pipe_198_inst RPIPE_ConvTranspose_input_pipe_286_inst RPIPE_ConvTranspose_input_pipe_299_inst RPIPE_ConvTranspose_input_pipe_311_inst RPIPE_ConvTranspose_input_pipe_324_inst RPIPE_ConvTranspose_input_pipe_336_inst RPIPE_ConvTranspose_input_pipe_349_inst RPIPE_ConvTranspose_input_pipe_361_inst RPIPE_ConvTranspose_input_pipe_374_inst RPIPE_ConvTranspose_input_pipe_386_inst RPIPE_ConvTranspose_input_pipe_399_inst 
    InportGroup_4: Block -- 
      signal data_out: std_logic_vector(319 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 39 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 39 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 39 downto 0);
      signal guard_vector : std_logic_vector( 39 downto 0);
      constant outBUFs : IntegerArray(39 downto 0) := (39 => 1, 38 => 1, 37 => 1, 36 => 1, 35 => 1, 34 => 1, 33 => 1, 32 => 1, 31 => 1, 30 => 1, 29 => 1, 28 => 1, 27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(39 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false, 28 => false, 29 => false, 30 => false, 31 => false, 32 => false, 33 => false, 34 => false, 35 => false, 36 => false, 37 => false, 38 => false, 39 => false);
      constant guardBuffering: IntegerArray(39 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2, 28 => 2, 29 => 2, 30 => 2, 31 => 2, 32 => 2, 33 => 2, 34 => 2, 35 => 2, 36 => 2, 37 => 2, 38 => 2, 39 => 2);
      -- 
    begin -- 
      reqL_unguarded(39) <= RPIPE_ConvTranspose_input_pipe_724_inst_req_0;
      reqL_unguarded(38) <= RPIPE_ConvTranspose_input_pipe_589_inst_req_0;
      reqL_unguarded(37) <= RPIPE_ConvTranspose_input_pipe_517_inst_req_0;
      reqL_unguarded(36) <= RPIPE_ConvTranspose_input_pipe_607_inst_req_0;
      reqL_unguarded(35) <= RPIPE_ConvTranspose_input_pipe_110_inst_req_0;
      reqL_unguarded(34) <= RPIPE_ConvTranspose_input_pipe_73_inst_req_0;
      reqL_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_135_inst_req_0;
      reqL_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_98_inst_req_0;
      reqL_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_486_inst_req_0;
      reqL_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_571_inst_req_0;
      reqL_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_742_inst_req_0;
      reqL_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_123_inst_req_0;
      reqL_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_48_inst_req_0;
      reqL_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_814_inst_req_0;
      reqL_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_693_inst_req_0;
      reqL_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_60_inst_req_0;
      reqL_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_85_inst_req_0;
      reqL_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_760_inst_req_0;
      reqL_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_535_inst_req_0;
      reqL_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_778_inst_req_0;
      reqL_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_35_inst_req_0;
      reqL_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_499_inst_req_0;
      reqL_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_553_inst_req_0;
      reqL_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_706_inst_req_0;
      reqL_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_796_inst_req_0;
      reqL_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_148_inst_req_0;
      reqL_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_160_inst_req_0;
      reqL_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_173_inst_req_0;
      reqL_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_185_inst_req_0;
      reqL_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_198_inst_req_0;
      reqL_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_286_inst_req_0;
      reqL_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_299_inst_req_0;
      reqL_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_311_inst_req_0;
      reqL_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_324_inst_req_0;
      reqL_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_336_inst_req_0;
      reqL_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_349_inst_req_0;
      reqL_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_361_inst_req_0;
      reqL_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_374_inst_req_0;
      reqL_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_386_inst_req_0;
      reqL_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_399_inst_req_0;
      RPIPE_ConvTranspose_input_pipe_724_inst_ack_0 <= ackL_unguarded(39);
      RPIPE_ConvTranspose_input_pipe_589_inst_ack_0 <= ackL_unguarded(38);
      RPIPE_ConvTranspose_input_pipe_517_inst_ack_0 <= ackL_unguarded(37);
      RPIPE_ConvTranspose_input_pipe_607_inst_ack_0 <= ackL_unguarded(36);
      RPIPE_ConvTranspose_input_pipe_110_inst_ack_0 <= ackL_unguarded(35);
      RPIPE_ConvTranspose_input_pipe_73_inst_ack_0 <= ackL_unguarded(34);
      RPIPE_ConvTranspose_input_pipe_135_inst_ack_0 <= ackL_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_98_inst_ack_0 <= ackL_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_486_inst_ack_0 <= ackL_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_571_inst_ack_0 <= ackL_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_742_inst_ack_0 <= ackL_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_123_inst_ack_0 <= ackL_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_48_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_814_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_693_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_60_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_85_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_760_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_535_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_778_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_35_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_499_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_553_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_706_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_796_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_148_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_160_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_173_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_185_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_198_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_286_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_299_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_311_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_324_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_336_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_349_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_361_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_374_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_386_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_399_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(39) <= RPIPE_ConvTranspose_input_pipe_724_inst_req_1;
      reqR_unguarded(38) <= RPIPE_ConvTranspose_input_pipe_589_inst_req_1;
      reqR_unguarded(37) <= RPIPE_ConvTranspose_input_pipe_517_inst_req_1;
      reqR_unguarded(36) <= RPIPE_ConvTranspose_input_pipe_607_inst_req_1;
      reqR_unguarded(35) <= RPIPE_ConvTranspose_input_pipe_110_inst_req_1;
      reqR_unguarded(34) <= RPIPE_ConvTranspose_input_pipe_73_inst_req_1;
      reqR_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_135_inst_req_1;
      reqR_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_98_inst_req_1;
      reqR_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_486_inst_req_1;
      reqR_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_571_inst_req_1;
      reqR_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_742_inst_req_1;
      reqR_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_123_inst_req_1;
      reqR_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_48_inst_req_1;
      reqR_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_814_inst_req_1;
      reqR_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_693_inst_req_1;
      reqR_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_60_inst_req_1;
      reqR_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_85_inst_req_1;
      reqR_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_760_inst_req_1;
      reqR_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_535_inst_req_1;
      reqR_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_778_inst_req_1;
      reqR_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_35_inst_req_1;
      reqR_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_499_inst_req_1;
      reqR_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_553_inst_req_1;
      reqR_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_706_inst_req_1;
      reqR_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_796_inst_req_1;
      reqR_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_148_inst_req_1;
      reqR_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_160_inst_req_1;
      reqR_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_173_inst_req_1;
      reqR_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_185_inst_req_1;
      reqR_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_198_inst_req_1;
      reqR_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_286_inst_req_1;
      reqR_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_299_inst_req_1;
      reqR_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_311_inst_req_1;
      reqR_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_324_inst_req_1;
      reqR_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_336_inst_req_1;
      reqR_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_349_inst_req_1;
      reqR_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_361_inst_req_1;
      reqR_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_374_inst_req_1;
      reqR_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_386_inst_req_1;
      reqR_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_399_inst_req_1;
      RPIPE_ConvTranspose_input_pipe_724_inst_ack_1 <= ackR_unguarded(39);
      RPIPE_ConvTranspose_input_pipe_589_inst_ack_1 <= ackR_unguarded(38);
      RPIPE_ConvTranspose_input_pipe_517_inst_ack_1 <= ackR_unguarded(37);
      RPIPE_ConvTranspose_input_pipe_607_inst_ack_1 <= ackR_unguarded(36);
      RPIPE_ConvTranspose_input_pipe_110_inst_ack_1 <= ackR_unguarded(35);
      RPIPE_ConvTranspose_input_pipe_73_inst_ack_1 <= ackR_unguarded(34);
      RPIPE_ConvTranspose_input_pipe_135_inst_ack_1 <= ackR_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_98_inst_ack_1 <= ackR_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_486_inst_ack_1 <= ackR_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_571_inst_ack_1 <= ackR_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_742_inst_ack_1 <= ackR_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_123_inst_ack_1 <= ackR_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_48_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_814_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_693_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_60_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_85_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_760_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_535_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_778_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_35_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_499_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_553_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_706_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_796_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_148_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_160_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_173_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_185_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_198_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_286_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_299_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_311_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_324_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_336_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_349_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_361_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_374_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_386_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_399_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      guard_vector(34)  <=  '1';
      guard_vector(35)  <=  '1';
      guard_vector(36)  <=  '1';
      guard_vector(37)  <=  '1';
      guard_vector(38)  <=  '1';
      guard_vector(39)  <=  '1';
      call209_725 <= data_out(319 downto 312);
      call177_590 <= data_out(311 downto 304);
      call153_518 <= data_out(303 downto 296);
      call183_608 <= data_out(295 downto 288);
      call23_111 <= data_out(287 downto 280);
      call10_74 <= data_out(279 downto 272);
      call32_136 <= data_out(271 downto 264);
      call19_99 <= data_out(263 downto 256);
      call143_487 <= data_out(255 downto 248);
      call171_572 <= data_out(247 downto 240);
      call215_743 <= data_out(239 downto 232);
      call28_124 <= data_out(231 downto 224);
      call2_49 <= data_out(223 downto 216);
      call239_815 <= data_out(215 downto 208);
      call199_694 <= data_out(207 downto 200);
      call5_61 <= data_out(199 downto 192);
      call14_86 <= data_out(191 downto 184);
      call221_761 <= data_out(183 downto 176);
      call159_536 <= data_out(175 downto 168);
      call227_779 <= data_out(167 downto 160);
      call_36 <= data_out(159 downto 152);
      call147_500 <= data_out(151 downto 144);
      call165_554 <= data_out(143 downto 136);
      call203_707 <= data_out(135 downto 128);
      call233_797 <= data_out(127 downto 120);
      call37_149 <= data_out(119 downto 112);
      call41_161 <= data_out(111 downto 104);
      call46_174 <= data_out(103 downto 96);
      call50_186 <= data_out(95 downto 88);
      call55_199 <= data_out(87 downto 80);
      call92_287 <= data_out(79 downto 72);
      call97_300 <= data_out(71 downto 64);
      call101_312 <= data_out(63 downto 56);
      call106_325 <= data_out(55 downto 48);
      call110_337 <= data_out(47 downto 40);
      call115_350 <= data_out(39 downto 32);
      call119_362 <= data_out(31 downto 24);
      call124_375 <= data_out(23 downto 16);
      call128_387 <= data_out(15 downto 8);
      call133_400 <= data_out(7 downto 0);
      ConvTranspose_input_pipe_read_4_gI: SplitGuardInterface generic map(name => "ConvTranspose_input_pipe_read_4_gI", nreqs => 40, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_input_pipe_read_4: InputPortRevised -- 
        generic map ( name => "ConvTranspose_input_pipe_read_4", data_width => 8,  num_reqs => 40,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => ConvTranspose_input_pipe_pipe_read_req(0),
          oack => ConvTranspose_input_pipe_pipe_read_ack(0),
          odata => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 4
    -- shared outport operator group (0) : WPIPE_Block0_start_995_inst WPIPE_Block0_start_998_inst WPIPE_Block0_start_1002_inst WPIPE_Block0_start_1006_inst WPIPE_Block0_start_971_inst WPIPE_Block0_start_1009_inst WPIPE_Block0_start_974_inst WPIPE_Block0_start_992_inst WPIPE_Block0_start_989_inst WPIPE_Block0_start_977_inst WPIPE_Block0_start_980_inst WPIPE_Block0_start_983_inst WPIPE_Block0_start_986_inst WPIPE_Block0_start_1012_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block0_start_995_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block0_start_998_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block0_start_1002_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block0_start_1006_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block0_start_971_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block0_start_1009_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block0_start_974_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block0_start_992_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block0_start_989_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block0_start_977_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block0_start_980_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block0_start_983_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block0_start_986_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block0_start_1012_inst_req_0;
      WPIPE_Block0_start_995_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block0_start_998_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block0_start_1002_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block0_start_1006_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block0_start_971_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block0_start_1009_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block0_start_974_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block0_start_992_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block0_start_989_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block0_start_977_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block0_start_980_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block0_start_983_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block0_start_986_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block0_start_1012_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block0_start_995_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block0_start_998_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block0_start_1002_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block0_start_1006_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block0_start_971_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block0_start_1009_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block0_start_974_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block0_start_992_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block0_start_989_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block0_start_977_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block0_start_980_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block0_start_983_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block0_start_986_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block0_start_1012_inst_req_1;
      WPIPE_Block0_start_995_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block0_start_998_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block0_start_1002_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block0_start_1006_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block0_start_971_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block0_start_1009_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block0_start_974_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block0_start_992_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block0_start_989_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block0_start_977_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block0_start_980_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block0_start_983_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block0_start_986_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block0_start_1012_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= add108_334 & type_cast_1000_wire_constant & type_cast_1004_wire_constant & add117_359 & add_58 & add126_384 & add12_83 & add99_309 & add57_208 & add21_108 & add30_133 & add39_158 & add48_183 & add135_409;
      Block0_start_write_0_gI: SplitGuardInterface generic map(name => "Block0_start_write_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_start_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_start_pipe_write_req(0),
          oack => Block0_start_pipe_write_ack(0),
          odata => Block0_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_Block1_start_1021_inst WPIPE_Block1_start_1024_inst WPIPE_Block1_start_1068_inst WPIPE_Block1_start_1033_inst WPIPE_Block1_start_1059_inst WPIPE_Block1_start_1027_inst WPIPE_Block1_start_1062_inst WPIPE_Block1_start_1036_inst WPIPE_Block1_start_1018_inst WPIPE_Block1_start_1039_inst WPIPE_Block1_start_1065_inst WPIPE_Block1_start_1030_inst WPIPE_Block1_start_1052_inst WPIPE_Block1_start_1015_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block1_start_1021_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block1_start_1024_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block1_start_1068_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block1_start_1033_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block1_start_1059_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block1_start_1027_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block1_start_1062_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block1_start_1036_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block1_start_1018_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block1_start_1039_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block1_start_1065_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block1_start_1030_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block1_start_1052_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block1_start_1015_inst_req_0;
      WPIPE_Block1_start_1021_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block1_start_1024_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block1_start_1068_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block1_start_1033_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block1_start_1059_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block1_start_1027_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block1_start_1062_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block1_start_1036_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block1_start_1018_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block1_start_1039_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block1_start_1065_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block1_start_1030_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block1_start_1052_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block1_start_1015_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block1_start_1021_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block1_start_1024_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block1_start_1068_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block1_start_1033_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block1_start_1059_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block1_start_1027_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block1_start_1062_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block1_start_1036_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block1_start_1018_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block1_start_1039_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block1_start_1065_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block1_start_1030_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block1_start_1052_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block1_start_1015_inst_req_1;
      WPIPE_Block1_start_1021_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block1_start_1024_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block1_start_1068_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block1_start_1033_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block1_start_1059_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block1_start_1027_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block1_start_1062_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block1_start_1036_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block1_start_1018_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block1_start_1039_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block1_start_1065_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block1_start_1030_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block1_start_1052_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block1_start_1015_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= add21_108 & add30_133 & add135_409 & add57_208 & conv307_1058 & add39_158 & add117_359 & add99_309 & add12_83 & add108_334 & add126_384 & add48_183 & conv305_1051 & add_58;
      Block1_start_write_1_gI: SplitGuardInterface generic map(name => "Block1_start_write_1_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_start_write_1: OutputPortRevised -- 
        generic map ( name => "Block1_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_start_pipe_write_req(0),
          oack => Block1_start_pipe_write_ack(0),
          odata => Block1_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_Block2_start_1115_inst WPIPE_Block2_start_1124_inst WPIPE_Block2_start_1086_inst WPIPE_Block2_start_1071_inst WPIPE_Block2_start_1080_inst WPIPE_Block2_start_1092_inst WPIPE_Block2_start_1077_inst WPIPE_Block2_start_1118_inst WPIPE_Block2_start_1095_inst WPIPE_Block2_start_1083_inst WPIPE_Block2_start_1089_inst WPIPE_Block2_start_1121_inst WPIPE_Block2_start_1074_inst WPIPE_Block2_start_1108_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block2_start_1115_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block2_start_1124_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block2_start_1086_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block2_start_1071_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block2_start_1080_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block2_start_1092_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block2_start_1077_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block2_start_1118_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block2_start_1095_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block2_start_1083_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block2_start_1089_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block2_start_1121_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block2_start_1074_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block2_start_1108_inst_req_0;
      WPIPE_Block2_start_1115_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block2_start_1124_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block2_start_1086_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block2_start_1071_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block2_start_1080_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block2_start_1092_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block2_start_1077_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block2_start_1118_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block2_start_1095_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block2_start_1083_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block2_start_1089_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block2_start_1121_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block2_start_1074_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block2_start_1108_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block2_start_1115_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block2_start_1124_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block2_start_1086_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block2_start_1071_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block2_start_1080_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block2_start_1092_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block2_start_1077_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block2_start_1118_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block2_start_1095_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block2_start_1083_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block2_start_1089_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block2_start_1121_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block2_start_1074_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block2_start_1108_inst_req_1;
      WPIPE_Block2_start_1115_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block2_start_1124_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block2_start_1086_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block2_start_1071_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block2_start_1080_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block2_start_1092_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block2_start_1077_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block2_start_1118_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block2_start_1095_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block2_start_1083_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block2_start_1089_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block2_start_1121_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block2_start_1074_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block2_start_1108_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= conv324_1114 & add135_409 & add48_183 & add_58 & add30_133 & add99_309 & add21_108 & add117_359 & add108_334 & add39_158 & add57_208 & add126_384 & add12_83 & conv322_1107;
      Block2_start_write_2_gI: SplitGuardInterface generic map(name => "Block2_start_write_2_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_start_write_2: OutputPortRevised -- 
        generic map ( name => "Block2_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_start_pipe_write_req(0),
          oack => Block2_start_pipe_write_ack(0),
          odata => Block2_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_Block3_start_1142_inst WPIPE_Block3_start_1127_inst WPIPE_Block3_start_1139_inst WPIPE_Block3_start_1151_inst WPIPE_Block3_start_1133_inst WPIPE_Block3_start_1130_inst WPIPE_Block3_start_1136_inst WPIPE_Block3_start_1180_inst WPIPE_Block3_start_1148_inst WPIPE_Block3_start_1145_inst WPIPE_Block3_start_1177_inst WPIPE_Block3_start_1174_inst WPIPE_Block3_start_1171_inst WPIPE_Block3_start_1164_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block3_start_1142_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block3_start_1127_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block3_start_1139_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block3_start_1151_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block3_start_1133_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block3_start_1130_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block3_start_1136_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block3_start_1180_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block3_start_1148_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block3_start_1145_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block3_start_1177_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block3_start_1174_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block3_start_1171_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block3_start_1164_inst_req_0;
      WPIPE_Block3_start_1142_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block3_start_1127_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block3_start_1139_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block3_start_1151_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block3_start_1133_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block3_start_1130_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block3_start_1136_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block3_start_1180_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block3_start_1148_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block3_start_1145_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block3_start_1177_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block3_start_1174_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block3_start_1171_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block3_start_1164_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block3_start_1142_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block3_start_1127_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block3_start_1139_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block3_start_1151_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block3_start_1133_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block3_start_1130_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block3_start_1136_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block3_start_1180_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block3_start_1148_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block3_start_1145_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block3_start_1177_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block3_start_1174_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block3_start_1171_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block3_start_1164_inst_req_1;
      WPIPE_Block3_start_1142_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block3_start_1127_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block3_start_1139_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block3_start_1151_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block3_start_1133_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block3_start_1130_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block3_start_1136_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block3_start_1180_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block3_start_1148_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block3_start_1145_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block3_start_1177_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block3_start_1174_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block3_start_1171_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block3_start_1164_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= add48_183 & add_58 & add39_158 & add108_334 & add21_108 & add12_83 & add30_133 & add135_409 & add99_309 & add57_208 & add126_384 & add117_359 & conv341_1170 & conv339_1163;
      Block3_start_write_3_gI: SplitGuardInterface generic map(name => "Block3_start_write_3_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_start_write_3: OutputPortRevised -- 
        generic map ( name => "Block3_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_start_pipe_write_req(0),
          oack => Block3_start_pipe_write_ack(0),
          odata => Block3_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared outport operator group (4) : WPIPE_ConvTranspose_output_pipe_1303_inst WPIPE_ConvTranspose_output_pipe_1300_inst WPIPE_ConvTranspose_output_pipe_1297_inst WPIPE_ConvTranspose_output_pipe_1294_inst WPIPE_ConvTranspose_output_pipe_1285_inst WPIPE_ConvTranspose_output_pipe_1291_inst WPIPE_ConvTranspose_output_pipe_1288_inst WPIPE_ConvTranspose_output_pipe_1306_inst WPIPE_ConvTranspose_output_pipe_1447_inst WPIPE_ConvTranspose_output_pipe_1450_inst WPIPE_ConvTranspose_output_pipe_1453_inst WPIPE_ConvTranspose_output_pipe_1456_inst WPIPE_ConvTranspose_output_pipe_1459_inst WPIPE_ConvTranspose_output_pipe_1462_inst WPIPE_ConvTranspose_output_pipe_1465_inst WPIPE_ConvTranspose_output_pipe_1468_inst 
    OutportGroup_4: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal sample_req, sample_ack : BooleanArray( 15 downto 0);
      signal update_req, update_ack : BooleanArray( 15 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 15 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 15 downto 0);
      signal guard_vector : std_logic_vector( 15 downto 0);
      constant inBUFs : IntegerArray(15 downto 0) := (15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(15 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false);
      constant guardBuffering: IntegerArray(15 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2);
      -- 
    begin -- 
      sample_req_unguarded(15) <= WPIPE_ConvTranspose_output_pipe_1303_inst_req_0;
      sample_req_unguarded(14) <= WPIPE_ConvTranspose_output_pipe_1300_inst_req_0;
      sample_req_unguarded(13) <= WPIPE_ConvTranspose_output_pipe_1297_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_ConvTranspose_output_pipe_1294_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_ConvTranspose_output_pipe_1285_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_ConvTranspose_output_pipe_1291_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_ConvTranspose_output_pipe_1288_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_ConvTranspose_output_pipe_1306_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1447_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1450_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1453_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1456_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1459_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1462_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1465_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1468_inst_req_0;
      WPIPE_ConvTranspose_output_pipe_1303_inst_ack_0 <= sample_ack_unguarded(15);
      WPIPE_ConvTranspose_output_pipe_1300_inst_ack_0 <= sample_ack_unguarded(14);
      WPIPE_ConvTranspose_output_pipe_1297_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_ConvTranspose_output_pipe_1294_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_ConvTranspose_output_pipe_1285_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_ConvTranspose_output_pipe_1291_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_ConvTranspose_output_pipe_1288_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_ConvTranspose_output_pipe_1306_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_ConvTranspose_output_pipe_1447_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1450_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1453_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1456_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1459_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1462_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1465_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1468_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(15) <= WPIPE_ConvTranspose_output_pipe_1303_inst_req_1;
      update_req_unguarded(14) <= WPIPE_ConvTranspose_output_pipe_1300_inst_req_1;
      update_req_unguarded(13) <= WPIPE_ConvTranspose_output_pipe_1297_inst_req_1;
      update_req_unguarded(12) <= WPIPE_ConvTranspose_output_pipe_1294_inst_req_1;
      update_req_unguarded(11) <= WPIPE_ConvTranspose_output_pipe_1285_inst_req_1;
      update_req_unguarded(10) <= WPIPE_ConvTranspose_output_pipe_1291_inst_req_1;
      update_req_unguarded(9) <= WPIPE_ConvTranspose_output_pipe_1288_inst_req_1;
      update_req_unguarded(8) <= WPIPE_ConvTranspose_output_pipe_1306_inst_req_1;
      update_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1447_inst_req_1;
      update_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1450_inst_req_1;
      update_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1453_inst_req_1;
      update_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1456_inst_req_1;
      update_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1459_inst_req_1;
      update_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1462_inst_req_1;
      update_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1465_inst_req_1;
      update_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1468_inst_req_1;
      WPIPE_ConvTranspose_output_pipe_1303_inst_ack_1 <= update_ack_unguarded(15);
      WPIPE_ConvTranspose_output_pipe_1300_inst_ack_1 <= update_ack_unguarded(14);
      WPIPE_ConvTranspose_output_pipe_1297_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_ConvTranspose_output_pipe_1294_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_ConvTranspose_output_pipe_1285_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_ConvTranspose_output_pipe_1291_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_ConvTranspose_output_pipe_1288_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_ConvTranspose_output_pipe_1306_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_ConvTranspose_output_pipe_1447_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1450_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1453_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1456_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1459_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1462_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1465_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1468_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      data_in <= conv368_1224 & conv374_1234 & conv380_1244 & conv386_1254 & conv404_1284 & conv392_1264 & conv398_1274 & conv362_1214 & conv480_1446 & conv474_1436 & conv468_1426 & conv462_1416 & conv456_1406 & conv450_1396 & conv444_1386 & conv438_1376;
      ConvTranspose_output_pipe_write_4_gI: SplitGuardInterface generic map(name => "ConvTranspose_output_pipe_write_4_gI", nreqs => 16, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_output_pipe_write_4: OutputPortRevised -- 
        generic map ( name => "ConvTranspose_output_pipe", data_width => 8, num_reqs => 16, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => ConvTranspose_output_pipe_pipe_write_req(0),
          oack => ConvTranspose_output_pipe_pipe_write_ack(0),
          odata => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 4
    -- shared outport operator group (5) : WPIPE_elapsed_time_pipe_1208_inst 
    OutportGroup_5: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1208_inst_req_0;
      WPIPE_elapsed_time_pipe_1208_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1208_inst_req_1;
      WPIPE_elapsed_time_pipe_1208_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= sub_1207;
      elapsed_time_pipe_write_5_gI: SplitGuardInterface generic map(name => "elapsed_time_pipe_write_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      elapsed_time_pipe_write_5: OutputPortRevised -- 
        generic map ( name => "elapsed_time_pipe", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => elapsed_time_pipe_pipe_write_req(0),
          oack => elapsed_time_pipe_pipe_write_ack(0),
          odata => elapsed_time_pipe_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 5
    -- shared call operator group (0) : call_stmt_963_call call_stmt_1197_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_963_call_req_0;
      reqL_unguarded(0) <= call_stmt_1197_call_req_0;
      call_stmt_963_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1197_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_963_call_req_1;
      reqR_unguarded(0) <= call_stmt_1197_call_req_1;
      call_stmt_963_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1197_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call275_963 <= data_out(127 downto 64);
      call354_1197 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end convTranspose_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeA is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeA;
architecture convTransposeA_arch of convTransposeA is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeA_CP_3777_start: Boolean;
  signal convTransposeA_CP_3777_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_1542_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1519_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1538_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1513_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1501_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1538_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1513_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1522_inst_req_0 : boolean;
  signal WPIPE_Block0_done_1843_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1522_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1522_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1550_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1553_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1553_inst_req_1 : boolean;
  signal type_cast_1542_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1550_inst_req_0 : boolean;
  signal type_cast_1632_inst_req_0 : boolean;
  signal phi_stmt_1612_ack_0 : boolean;
  signal type_cast_1820_inst_ack_0 : boolean;
  signal type_cast_1529_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1510_inst_ack_0 : boolean;
  signal type_cast_1632_inst_ack_0 : boolean;
  signal phi_stmt_1605_ack_0 : boolean;
  signal RPIPE_Block0_start_1519_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1510_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1522_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1507_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1507_inst_req_1 : boolean;
  signal type_cast_1830_inst_ack_1 : boolean;
  signal WPIPE_Block0_done_1843_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1510_inst_req_1 : boolean;
  signal phi_stmt_1626_req_0 : boolean;
  signal type_cast_1542_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1510_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1513_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1504_inst_ack_1 : boolean;
  signal type_cast_1632_inst_req_1 : boolean;
  signal phi_stmt_1626_ack_0 : boolean;
  signal type_cast_1611_inst_ack_1 : boolean;
  signal phi_stmt_1619_ack_0 : boolean;
  signal type_cast_1830_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1519_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1525_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1501_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1525_inst_ack_0 : boolean;
  signal type_cast_1529_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1498_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1519_inst_ack_1 : boolean;
  signal type_cast_1583_inst_ack_1 : boolean;
  signal type_cast_1583_inst_req_1 : boolean;
  signal type_cast_1529_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1498_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1550_inst_req_1 : boolean;
  signal type_cast_1583_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1550_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1516_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1501_inst_req_0 : boolean;
  signal type_cast_1529_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1516_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1556_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1516_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1504_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1513_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1504_inst_ack_0 : boolean;
  signal type_cast_1542_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1556_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1525_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1516_inst_ack_1 : boolean;
  signal type_cast_1832_inst_req_1 : boolean;
  signal type_cast_1583_inst_req_0 : boolean;
  signal type_cast_1820_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1556_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1538_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1507_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1525_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1498_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1538_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1504_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1501_inst_ack_0 : boolean;
  signal type_cast_1611_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1553_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1507_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1553_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1556_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1498_inst_ack_1 : boolean;
  signal type_cast_1820_inst_req_1 : boolean;
  signal phi_stmt_1605_req_0 : boolean;
  signal phi_stmt_1612_req_0 : boolean;
  signal type_cast_1820_inst_ack_1 : boolean;
  signal phi_stmt_1814_req_1 : boolean;
  signal phi_stmt_1827_req_0 : boolean;
  signal phi_stmt_1821_req_0 : boolean;
  signal type_cast_1587_inst_req_0 : boolean;
  signal type_cast_1587_inst_ack_0 : boolean;
  signal type_cast_1824_inst_ack_1 : boolean;
  signal type_cast_1587_inst_req_1 : boolean;
  signal type_cast_1830_inst_ack_0 : boolean;
  signal type_cast_1587_inst_ack_1 : boolean;
  signal type_cast_1824_inst_req_1 : boolean;
  signal type_cast_1591_inst_req_0 : boolean;
  signal type_cast_1830_inst_req_0 : boolean;
  signal type_cast_1591_inst_ack_0 : boolean;
  signal type_cast_1591_inst_req_1 : boolean;
  signal type_cast_1591_inst_ack_1 : boolean;
  signal phi_stmt_1814_req_0 : boolean;
  signal type_cast_1595_inst_req_0 : boolean;
  signal type_cast_1595_inst_ack_0 : boolean;
  signal type_cast_1824_inst_ack_0 : boolean;
  signal type_cast_1595_inst_req_1 : boolean;
  signal type_cast_1595_inst_ack_1 : boolean;
  signal type_cast_1832_inst_ack_0 : boolean;
  signal type_cast_1824_inst_req_0 : boolean;
  signal type_cast_1667_inst_req_0 : boolean;
  signal type_cast_1667_inst_ack_0 : boolean;
  signal type_cast_1667_inst_req_1 : boolean;
  signal type_cast_1667_inst_ack_1 : boolean;
  signal type_cast_1671_inst_req_0 : boolean;
  signal type_cast_1671_inst_ack_0 : boolean;
  signal type_cast_1671_inst_req_1 : boolean;
  signal type_cast_1671_inst_ack_1 : boolean;
  signal phi_stmt_1821_req_1 : boolean;
  signal type_cast_1826_inst_ack_1 : boolean;
  signal type_cast_1826_inst_req_1 : boolean;
  signal type_cast_1675_inst_req_0 : boolean;
  signal type_cast_1675_inst_ack_0 : boolean;
  signal type_cast_1675_inst_req_1 : boolean;
  signal type_cast_1675_inst_ack_1 : boolean;
  signal type_cast_1826_inst_ack_0 : boolean;
  signal type_cast_1705_inst_req_0 : boolean;
  signal type_cast_1705_inst_ack_0 : boolean;
  signal type_cast_1705_inst_req_1 : boolean;
  signal type_cast_1705_inst_ack_1 : boolean;
  signal phi_stmt_1827_ack_0 : boolean;
  signal phi_stmt_1821_ack_0 : boolean;
  signal type_cast_1826_inst_req_0 : boolean;
  signal phi_stmt_1619_req_1 : boolean;
  signal phi_stmt_1626_req_1 : boolean;
  signal type_cast_1625_inst_ack_1 : boolean;
  signal type_cast_1632_inst_ack_1 : boolean;
  signal type_cast_1625_inst_req_1 : boolean;
  signal array_obj_ref_1711_index_offset_req_0 : boolean;
  signal array_obj_ref_1711_index_offset_ack_0 : boolean;
  signal phi_stmt_1619_req_0 : boolean;
  signal array_obj_ref_1711_index_offset_req_1 : boolean;
  signal array_obj_ref_1711_index_offset_ack_1 : boolean;
  signal type_cast_1832_inst_req_0 : boolean;
  signal addr_of_1712_final_reg_req_0 : boolean;
  signal addr_of_1712_final_reg_ack_0 : boolean;
  signal phi_stmt_1827_req_1 : boolean;
  signal addr_of_1712_final_reg_req_1 : boolean;
  signal addr_of_1712_final_reg_ack_1 : boolean;
  signal phi_stmt_1814_ack_0 : boolean;
  signal type_cast_1625_inst_ack_0 : boolean;
  signal type_cast_1625_inst_req_0 : boolean;
  signal type_cast_1611_inst_ack_0 : boolean;
  signal ptr_deref_1716_load_0_req_0 : boolean;
  signal phi_stmt_1612_req_1 : boolean;
  signal ptr_deref_1716_load_0_ack_0 : boolean;
  signal WPIPE_Block0_done_1843_inst_ack_0 : boolean;
  signal type_cast_1611_inst_req_0 : boolean;
  signal ptr_deref_1716_load_0_req_1 : boolean;
  signal type_cast_1618_inst_ack_1 : boolean;
  signal ptr_deref_1716_load_0_ack_1 : boolean;
  signal type_cast_1832_inst_ack_1 : boolean;
  signal type_cast_1618_inst_req_1 : boolean;
  signal WPIPE_Block0_done_1843_inst_req_0 : boolean;
  signal type_cast_1618_inst_ack_0 : boolean;
  signal type_cast_1618_inst_req_0 : boolean;
  signal phi_stmt_1605_req_1 : boolean;
  signal array_obj_ref_1734_index_offset_req_0 : boolean;
  signal array_obj_ref_1734_index_offset_ack_0 : boolean;
  signal array_obj_ref_1734_index_offset_req_1 : boolean;
  signal array_obj_ref_1734_index_offset_ack_1 : boolean;
  signal addr_of_1735_final_reg_req_0 : boolean;
  signal addr_of_1735_final_reg_ack_0 : boolean;
  signal addr_of_1735_final_reg_req_1 : boolean;
  signal addr_of_1735_final_reg_ack_1 : boolean;
  signal ptr_deref_1738_store_0_req_0 : boolean;
  signal ptr_deref_1738_store_0_ack_0 : boolean;
  signal ptr_deref_1738_store_0_req_1 : boolean;
  signal ptr_deref_1738_store_0_ack_1 : boolean;
  signal type_cast_1743_inst_req_0 : boolean;
  signal type_cast_1743_inst_ack_0 : boolean;
  signal type_cast_1743_inst_req_1 : boolean;
  signal type_cast_1743_inst_ack_1 : boolean;
  signal if_stmt_1756_branch_req_0 : boolean;
  signal if_stmt_1756_branch_ack_1 : boolean;
  signal if_stmt_1756_branch_ack_0 : boolean;
  signal type_cast_1784_inst_req_0 : boolean;
  signal type_cast_1784_inst_ack_0 : boolean;
  signal type_cast_1784_inst_req_1 : boolean;
  signal type_cast_1784_inst_ack_1 : boolean;
  signal type_cast_1800_inst_req_0 : boolean;
  signal type_cast_1800_inst_ack_0 : boolean;
  signal type_cast_1800_inst_req_1 : boolean;
  signal type_cast_1800_inst_ack_1 : boolean;
  signal if_stmt_1807_branch_req_0 : boolean;
  signal if_stmt_1807_branch_ack_1 : boolean;
  signal if_stmt_1807_branch_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeA_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeA_CP_3777_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeA_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_3777_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeA_CP_3777_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_3777_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeA_CP_3777: Block -- control-path 
    signal convTransposeA_CP_3777_elements: BooleanArray(125 downto 0);
    -- 
  begin -- 
    convTransposeA_CP_3777_elements(0) <= convTransposeA_CP_3777_start;
    convTransposeA_CP_3777_symbol <= convTransposeA_CP_3777_elements(78);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/$entry
      -- CP-element group 0: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1498_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557__entry__
      -- CP-element group 0: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1498_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/type_cast_1542_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/type_cast_1542_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1496/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1496/branch_block_stmt_1496__entry__
      -- CP-element group 0: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/type_cast_1542_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1498_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/type_cast_1529_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/type_cast_1529_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/type_cast_1529_update_start_
      -- 
    cr_3998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(0), ack => type_cast_1542_inst_req_1); -- 
    rr_3825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(0), ack => RPIPE_Block0_start_1498_inst_req_0); -- 
    cr_3970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(0), ack => type_cast_1529_inst_req_1); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	125 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	84 
    -- CP-element group 1: 	85 
    -- CP-element group 1: 	87 
    -- CP-element group 1: 	88 
    -- CP-element group 1: 	90 
    -- CP-element group 1: 	91 
    -- CP-element group 1: 	93 
    -- CP-element group 1: 	94 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1626/phi_stmt_1626_sources/type_cast_1632/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1626/phi_stmt_1626_sources/type_cast_1632/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1626/phi_stmt_1626_sources/type_cast_1632/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1626/phi_stmt_1626_sources/type_cast_1632/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1605/$entry
      -- CP-element group 1: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1605/phi_stmt_1605_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1605/phi_stmt_1605_sources/type_cast_1611/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1496/merge_stmt_1813__exit__
      -- CP-element group 1: 	 branch_block_stmt_1496/assign_stmt_1839__entry__
      -- CP-element group 1: 	 branch_block_stmt_1496/assign_stmt_1839__exit__
      -- CP-element group 1: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1605/phi_stmt_1605_sources/type_cast_1611/$entry
      -- CP-element group 1: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1605/phi_stmt_1605_sources/type_cast_1611/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1605/phi_stmt_1605_sources/type_cast_1611/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1626/phi_stmt_1626_sources/type_cast_1632/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1626/phi_stmt_1626_sources/type_cast_1632/$entry
      -- CP-element group 1: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1626/phi_stmt_1626_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1626/$entry
      -- CP-element group 1: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1619/phi_stmt_1619_sources/type_cast_1625/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1619/phi_stmt_1619_sources/type_cast_1625/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1619/phi_stmt_1619_sources/type_cast_1625/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1619/phi_stmt_1619_sources/type_cast_1625/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1619/phi_stmt_1619_sources/type_cast_1625/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1619/phi_stmt_1619_sources/type_cast_1625/$entry
      -- CP-element group 1: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1619/phi_stmt_1619_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1619/$entry
      -- CP-element group 1: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1605/phi_stmt_1605_sources/type_cast_1611/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1605/phi_stmt_1605_sources/type_cast_1611/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1612/phi_stmt_1612_sources/type_cast_1618/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1612/phi_stmt_1612_sources/type_cast_1618/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1612/phi_stmt_1612_sources/type_cast_1618/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1612/phi_stmt_1612_sources/type_cast_1618/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1612/phi_stmt_1612_sources/type_cast_1618/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1612/phi_stmt_1612_sources/type_cast_1618/$entry
      -- CP-element group 1: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1612/phi_stmt_1612_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1612/$entry
      -- CP-element group 1: 	 branch_block_stmt_1496/assign_stmt_1839/$entry
      -- CP-element group 1: 	 branch_block_stmt_1496/assign_stmt_1839/$exit
      -- 
    rr_4580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(1), ack => type_cast_1632_inst_req_0); -- 
    cr_4585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(1), ack => type_cast_1632_inst_req_1); -- 
    cr_4516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(1), ack => type_cast_1611_inst_req_1); -- 
    cr_4562_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4562_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(1), ack => type_cast_1625_inst_req_1); -- 
    rr_4557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(1), ack => type_cast_1625_inst_req_0); -- 
    rr_4511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(1), ack => type_cast_1611_inst_req_0); -- 
    cr_4539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(1), ack => type_cast_1618_inst_req_1); -- 
    rr_4534_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4534_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(1), ack => type_cast_1618_inst_req_0); -- 
    convTransposeA_CP_3777_elements(1) <= convTransposeA_CP_3777_elements(125);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1498_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1498_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1498_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1498_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1498_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1498_Update/cr
      -- 
    ra_3826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1498_inst_ack_0, ack => convTransposeA_CP_3777_elements(2)); -- 
    cr_3830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(2), ack => RPIPE_Block0_start_1498_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1498_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1501_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1501_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1501_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1498_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1498_Update/ca
      -- 
    ca_3831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1498_inst_ack_1, ack => convTransposeA_CP_3777_elements(3)); -- 
    rr_3839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(3), ack => RPIPE_Block0_start_1501_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1501_update_start_
      -- CP-element group 4: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1501_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1501_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1501_Update/cr
      -- CP-element group 4: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1501_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1501_Update/$entry
      -- 
    ra_3840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1501_inst_ack_0, ack => convTransposeA_CP_3777_elements(4)); -- 
    cr_3844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(4), ack => RPIPE_Block0_start_1501_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1501_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1501_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1504_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1501_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1504_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1504_Sample/rr
      -- 
    ca_3845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1501_inst_ack_1, ack => convTransposeA_CP_3777_elements(5)); -- 
    rr_3853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(5), ack => RPIPE_Block0_start_1504_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1504_update_start_
      -- CP-element group 6: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1504_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1504_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1504_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1504_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1504_Update/cr
      -- 
    ra_3854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1504_inst_ack_0, ack => convTransposeA_CP_3777_elements(6)); -- 
    cr_3858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(6), ack => RPIPE_Block0_start_1504_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1507_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1504_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1504_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1507_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1504_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1507_Sample/rr
      -- 
    ca_3859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1504_inst_ack_1, ack => convTransposeA_CP_3777_elements(7)); -- 
    rr_3867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(7), ack => RPIPE_Block0_start_1507_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1507_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1507_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1507_Update/cr
      -- CP-element group 8: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1507_update_start_
      -- CP-element group 8: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1507_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1507_Sample/ra
      -- 
    ra_3868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1507_inst_ack_0, ack => convTransposeA_CP_3777_elements(8)); -- 
    cr_3872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(8), ack => RPIPE_Block0_start_1507_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1510_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1510_Sample/rr
      -- CP-element group 9: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1507_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1510_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1507_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1507_update_completed_
      -- 
    ca_3873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1507_inst_ack_1, ack => convTransposeA_CP_3777_elements(9)); -- 
    rr_3881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(9), ack => RPIPE_Block0_start_1510_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1510_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1510_update_start_
      -- CP-element group 10: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1510_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1510_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1510_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1510_Update/cr
      -- 
    ra_3882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1510_inst_ack_0, ack => convTransposeA_CP_3777_elements(10)); -- 
    cr_3886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(10), ack => RPIPE_Block0_start_1510_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1510_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1510_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1510_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1513_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1513_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1513_Sample/rr
      -- 
    ca_3887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1510_inst_ack_1, ack => convTransposeA_CP_3777_elements(11)); -- 
    rr_3895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(11), ack => RPIPE_Block0_start_1513_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1513_Update/cr
      -- CP-element group 12: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1513_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1513_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1513_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1513_update_start_
      -- CP-element group 12: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1513_Sample/$exit
      -- 
    ra_3896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1513_inst_ack_0, ack => convTransposeA_CP_3777_elements(12)); -- 
    cr_3900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(12), ack => RPIPE_Block0_start_1513_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1513_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1516_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1513_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1516_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1513_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1516_Sample/rr
      -- 
    ca_3901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1513_inst_ack_1, ack => convTransposeA_CP_3777_elements(13)); -- 
    rr_3909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(13), ack => RPIPE_Block0_start_1516_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1516_update_start_
      -- CP-element group 14: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1516_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1516_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1516_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1516_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1516_Update/cr
      -- 
    ra_3910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1516_inst_ack_0, ack => convTransposeA_CP_3777_elements(14)); -- 
    cr_3914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(14), ack => RPIPE_Block0_start_1516_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1519_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1516_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1516_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1516_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1519_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1519_Sample/$entry
      -- 
    ca_3915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1516_inst_ack_1, ack => convTransposeA_CP_3777_elements(15)); -- 
    rr_3923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(15), ack => RPIPE_Block0_start_1519_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1519_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1519_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1519_Update/cr
      -- CP-element group 16: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1519_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1519_update_start_
      -- CP-element group 16: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1519_Sample/$exit
      -- 
    ra_3924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1519_inst_ack_0, ack => convTransposeA_CP_3777_elements(16)); -- 
    cr_3928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(16), ack => RPIPE_Block0_start_1519_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1522_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1519_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1519_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1522_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1522_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1519_update_completed_
      -- 
    ca_3929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1519_inst_ack_1, ack => convTransposeA_CP_3777_elements(17)); -- 
    rr_3937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(17), ack => RPIPE_Block0_start_1522_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1522_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1522_Update/cr
      -- CP-element group 18: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1522_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1522_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1522_update_start_
      -- CP-element group 18: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1522_Sample/$exit
      -- 
    ra_3938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1522_inst_ack_0, ack => convTransposeA_CP_3777_elements(18)); -- 
    cr_3942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(18), ack => RPIPE_Block0_start_1522_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1525_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1522_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1525_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1525_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1522_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1522_update_completed_
      -- 
    ca_3943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1522_inst_ack_1, ack => convTransposeA_CP_3777_elements(19)); -- 
    rr_3951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(19), ack => RPIPE_Block0_start_1525_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1525_update_start_
      -- CP-element group 20: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1525_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1525_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1525_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1525_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1525_Update/cr
      -- 
    ra_3952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1525_inst_ack_0, ack => convTransposeA_CP_3777_elements(20)); -- 
    cr_3956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(20), ack => RPIPE_Block0_start_1525_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/type_cast_1529_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1525_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1525_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1538_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1538_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1538_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1525_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/type_cast_1529_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/type_cast_1529_Sample/$entry
      -- 
    ca_3957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1525_inst_ack_1, ack => convTransposeA_CP_3777_elements(21)); -- 
    rr_3965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(21), ack => type_cast_1529_inst_req_0); -- 
    rr_3979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(21), ack => RPIPE_Block0_start_1538_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/type_cast_1529_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/type_cast_1529_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/type_cast_1529_sample_completed_
      -- 
    ra_3966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1529_inst_ack_0, ack => convTransposeA_CP_3777_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/type_cast_1529_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/type_cast_1529_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/type_cast_1529_update_completed_
      -- 
    ca_3971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1529_inst_ack_1, ack => convTransposeA_CP_3777_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1538_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1538_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1538_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1538_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1538_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1538_Sample/ra
      -- 
    ra_3980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1538_inst_ack_0, ack => convTransposeA_CP_3777_elements(24)); -- 
    cr_3984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(24), ack => RPIPE_Block0_start_1538_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1550_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1550_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1538_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1550_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/type_cast_1542_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1538_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/type_cast_1542_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/type_cast_1542_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1538_update_completed_
      -- 
    ca_3985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1538_inst_ack_1, ack => convTransposeA_CP_3777_elements(25)); -- 
    rr_3993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(25), ack => type_cast_1542_inst_req_0); -- 
    rr_4007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(25), ack => RPIPE_Block0_start_1550_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/type_cast_1542_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/type_cast_1542_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/type_cast_1542_Sample/ra
      -- 
    ra_3994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1542_inst_ack_0, ack => convTransposeA_CP_3777_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/type_cast_1542_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/type_cast_1542_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/type_cast_1542_Update/$exit
      -- 
    ca_3999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1542_inst_ack_1, ack => convTransposeA_CP_3777_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1550_update_start_
      -- CP-element group 28: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1550_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1550_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1550_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1550_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1550_Update/cr
      -- 
    ra_4008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1550_inst_ack_0, ack => convTransposeA_CP_3777_elements(28)); -- 
    cr_4012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(28), ack => RPIPE_Block0_start_1550_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1550_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1550_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1550_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1553_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1553_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1553_Sample/rr
      -- 
    ca_4013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1550_inst_ack_1, ack => convTransposeA_CP_3777_elements(29)); -- 
    rr_4021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(29), ack => RPIPE_Block0_start_1553_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1553_Update/cr
      -- CP-element group 30: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1553_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1553_update_start_
      -- CP-element group 30: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1553_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1553_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1553_Update/$entry
      -- 
    ra_4022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1553_inst_ack_0, ack => convTransposeA_CP_3777_elements(30)); -- 
    cr_4026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(30), ack => RPIPE_Block0_start_1553_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1553_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1556_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1553_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1556_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1556_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1553_update_completed_
      -- 
    ca_4027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1553_inst_ack_1, ack => convTransposeA_CP_3777_elements(31)); -- 
    rr_4035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(31), ack => RPIPE_Block0_start_1556_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1556_update_start_
      -- CP-element group 32: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1556_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1556_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1556_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1556_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1556_Update/cr
      -- 
    ra_4036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1556_inst_ack_0, ack => convTransposeA_CP_3777_elements(32)); -- 
    cr_4040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(32), ack => RPIPE_Block0_start_1556_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1556_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1556_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/RPIPE_Block0_start_1556_Update/$exit
      -- 
    ca_4041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1556_inst_ack_1, ack => convTransposeA_CP_3777_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34: 	41 
    -- CP-element group 34: 	42 
    -- CP-element group 34:  members (28) 
      -- CP-element group 34: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557/$exit
      -- CP-element group 34: 	 branch_block_stmt_1496/assign_stmt_1499_to_assign_stmt_1557__exit__
      -- CP-element group 34: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602__entry__
      -- CP-element group 34: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1583_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1583_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1583_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1583_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1583_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/$entry
      -- CP-element group 34: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1583_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1587_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1587_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1587_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1587_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1587_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1587_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1591_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1591_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1591_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1591_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1591_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1591_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1595_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1595_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1595_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1595_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1595_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1595_Update/cr
      -- 
    cr_4057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(34), ack => type_cast_1583_inst_req_1); -- 
    rr_4052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(34), ack => type_cast_1583_inst_req_0); -- 
    rr_4066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(34), ack => type_cast_1587_inst_req_0); -- 
    cr_4071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(34), ack => type_cast_1587_inst_req_1); -- 
    rr_4080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(34), ack => type_cast_1591_inst_req_0); -- 
    cr_4085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(34), ack => type_cast_1591_inst_req_1); -- 
    rr_4094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(34), ack => type_cast_1595_inst_req_0); -- 
    cr_4099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(34), ack => type_cast_1595_inst_req_1); -- 
    convTransposeA_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3777_elements(23) & convTransposeA_CP_3777_elements(27) & convTransposeA_CP_3777_elements(33);
      gj_convTransposeA_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3777_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1583_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1583_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1583_Sample/$exit
      -- 
    ra_4053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1583_inst_ack_0, ack => convTransposeA_CP_3777_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	43 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1583_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1583_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1583_update_completed_
      -- 
    ca_4058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1583_inst_ack_1, ack => convTransposeA_CP_3777_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1587_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1587_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1587_Sample/ra
      -- 
    ra_4067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1587_inst_ack_0, ack => convTransposeA_CP_3777_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	43 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1587_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1587_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1587_Update/ca
      -- 
    ca_4072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1587_inst_ack_1, ack => convTransposeA_CP_3777_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1591_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1591_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1591_Sample/ra
      -- 
    ra_4081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1591_inst_ack_0, ack => convTransposeA_CP_3777_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	43 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1591_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1591_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1591_Update/ca
      -- 
    ca_4086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1591_inst_ack_1, ack => convTransposeA_CP_3777_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	34 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1595_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1595_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1595_Sample/ra
      -- 
    ra_4095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1595_inst_ack_0, ack => convTransposeA_CP_3777_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	34 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1595_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1595_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/type_cast_1595_Update/ca
      -- 
    ca_4100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1595_inst_ack_1, ack => convTransposeA_CP_3777_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  place  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	36 
    -- CP-element group 43: 	38 
    -- CP-element group 43: 	40 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	79 
    -- CP-element group 43: 	80 
    -- CP-element group 43: 	81 
    -- CP-element group 43: 	82 
    -- CP-element group 43:  members (12) 
      -- CP-element group 43: 	 branch_block_stmt_1496/entry_whilex_xbody
      -- CP-element group 43: 	 branch_block_stmt_1496/entry_whilex_xbody_PhiReq/phi_stmt_1605/phi_stmt_1605_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1496/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 43: 	 branch_block_stmt_1496/entry_whilex_xbody_PhiReq/phi_stmt_1605/$entry
      -- CP-element group 43: 	 branch_block_stmt_1496/entry_whilex_xbody_PhiReq/phi_stmt_1612/phi_stmt_1612_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1496/entry_whilex_xbody_PhiReq/phi_stmt_1626/phi_stmt_1626_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602__exit__
      -- CP-element group 43: 	 branch_block_stmt_1496/assign_stmt_1564_to_assign_stmt_1602/$exit
      -- CP-element group 43: 	 branch_block_stmt_1496/entry_whilex_xbody_PhiReq/phi_stmt_1612/$entry
      -- CP-element group 43: 	 branch_block_stmt_1496/entry_whilex_xbody_PhiReq/phi_stmt_1626/$entry
      -- CP-element group 43: 	 branch_block_stmt_1496/entry_whilex_xbody_PhiReq/phi_stmt_1619/phi_stmt_1619_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1496/entry_whilex_xbody_PhiReq/phi_stmt_1619/$entry
      -- 
    convTransposeA_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3777_elements(36) & convTransposeA_CP_3777_elements(38) & convTransposeA_CP_3777_elements(40) & convTransposeA_CP_3777_elements(42);
      gj_convTransposeA_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3777_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	102 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1667_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1667_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1667_Sample/ra
      -- 
    ra_4112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1667_inst_ack_0, ack => convTransposeA_CP_3777_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	102 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	58 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1667_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1667_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1667_Update/ca
      -- 
    ca_4117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1667_inst_ack_1, ack => convTransposeA_CP_3777_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	102 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1671_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1671_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1671_Sample/ra
      -- 
    ra_4126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1671_inst_ack_0, ack => convTransposeA_CP_3777_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	102 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	58 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1671_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1671_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1671_Update/ca
      -- 
    ca_4131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1671_inst_ack_1, ack => convTransposeA_CP_3777_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	102 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1675_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1675_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1675_Sample/ra
      -- 
    ra_4140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1675_inst_ack_0, ack => convTransposeA_CP_3777_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	102 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1675_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1675_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1675_Update/ca
      -- 
    ca_4145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1675_inst_ack_1, ack => convTransposeA_CP_3777_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	102 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1705_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1705_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1705_Sample/ra
      -- 
    ra_4154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1705_inst_ack_0, ack => convTransposeA_CP_3777_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	102 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (16) 
      -- CP-element group 51: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1705_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1705_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1705_Update/ca
      -- CP-element group 51: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1711_index_resized_1
      -- CP-element group 51: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1711_index_scaled_1
      -- CP-element group 51: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1711_index_computed_1
      -- CP-element group 51: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1711_index_resize_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1711_index_resize_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1711_index_resize_1/index_resize_req
      -- CP-element group 51: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1711_index_resize_1/index_resize_ack
      -- CP-element group 51: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1711_index_scale_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1711_index_scale_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1711_index_scale_1/scale_rename_req
      -- CP-element group 51: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1711_index_scale_1/scale_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1711_final_index_sum_regn_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1711_final_index_sum_regn_Sample/req
      -- 
    ca_4159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1705_inst_ack_1, ack => convTransposeA_CP_3777_elements(51)); -- 
    req_4184_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4184_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(51), ack => array_obj_ref_1711_index_offset_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	68 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1711_final_index_sum_regn_sample_complete
      -- CP-element group 52: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1711_final_index_sum_regn_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1711_final_index_sum_regn_Sample/ack
      -- 
    ack_4185_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1711_index_offset_ack_0, ack => convTransposeA_CP_3777_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	102 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (11) 
      -- CP-element group 53: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/addr_of_1712_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1711_root_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1711_offset_calculated
      -- CP-element group 53: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1711_final_index_sum_regn_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1711_final_index_sum_regn_Update/ack
      -- CP-element group 53: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1711_base_plus_offset/$entry
      -- CP-element group 53: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1711_base_plus_offset/$exit
      -- CP-element group 53: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1711_base_plus_offset/sum_rename_req
      -- CP-element group 53: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1711_base_plus_offset/sum_rename_ack
      -- CP-element group 53: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/addr_of_1712_request/$entry
      -- CP-element group 53: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/addr_of_1712_request/req
      -- 
    ack_4190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1711_index_offset_ack_1, ack => convTransposeA_CP_3777_elements(53)); -- 
    req_4199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(53), ack => addr_of_1712_final_reg_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/addr_of_1712_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/addr_of_1712_request/$exit
      -- CP-element group 54: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/addr_of_1712_request/ack
      -- 
    ack_4200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1712_final_reg_ack_0, ack => convTransposeA_CP_3777_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	102 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (24) 
      -- CP-element group 55: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/addr_of_1712_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/addr_of_1712_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/addr_of_1712_complete/ack
      -- CP-element group 55: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1716_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1716_base_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1716_word_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1716_root_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1716_base_address_resized
      -- CP-element group 55: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1716_base_addr_resize/$entry
      -- CP-element group 55: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1716_base_addr_resize/$exit
      -- CP-element group 55: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1716_base_addr_resize/base_resize_req
      -- CP-element group 55: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1716_base_addr_resize/base_resize_ack
      -- CP-element group 55: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1716_base_plus_offset/$entry
      -- CP-element group 55: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1716_base_plus_offset/$exit
      -- CP-element group 55: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1716_base_plus_offset/sum_rename_req
      -- CP-element group 55: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1716_base_plus_offset/sum_rename_ack
      -- CP-element group 55: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1716_word_addrgen/$entry
      -- CP-element group 55: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1716_word_addrgen/$exit
      -- CP-element group 55: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1716_word_addrgen/root_register_req
      -- CP-element group 55: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1716_word_addrgen/root_register_ack
      -- CP-element group 55: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1716_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1716_Sample/word_access_start/$entry
      -- CP-element group 55: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1716_Sample/word_access_start/word_0/$entry
      -- CP-element group 55: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1716_Sample/word_access_start/word_0/rr
      -- 
    ack_4205_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1712_final_reg_ack_1, ack => convTransposeA_CP_3777_elements(55)); -- 
    rr_4238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(55), ack => ptr_deref_1716_load_0_req_0); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (5) 
      -- CP-element group 56: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1716_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1716_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1716_Sample/word_access_start/$exit
      -- CP-element group 56: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1716_Sample/word_access_start/word_0/$exit
      -- CP-element group 56: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1716_Sample/word_access_start/word_0/ra
      -- 
    ra_4239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1716_load_0_ack_0, ack => convTransposeA_CP_3777_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	102 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (9) 
      -- CP-element group 57: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1716_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1716_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1716_Update/word_access_complete/$exit
      -- CP-element group 57: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1716_Update/word_access_complete/word_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1716_Update/word_access_complete/word_0/ca
      -- CP-element group 57: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1716_Update/ptr_deref_1716_Merge/$entry
      -- CP-element group 57: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1716_Update/ptr_deref_1716_Merge/$exit
      -- CP-element group 57: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1716_Update/ptr_deref_1716_Merge/merge_req
      -- CP-element group 57: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1716_Update/ptr_deref_1716_Merge/merge_ack
      -- 
    ca_4250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1716_load_0_ack_1, ack => convTransposeA_CP_3777_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	45 
    -- CP-element group 58: 	47 
    -- CP-element group 58: 	49 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (13) 
      -- CP-element group 58: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1734_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1734_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1734_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1734_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1734_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1734_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1734_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1734_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1734_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1734_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1734_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1734_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1734_final_index_sum_regn_Sample/req
      -- 
    req_4280_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4280_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(58), ack => array_obj_ref_1734_index_offset_req_0); -- 
    convTransposeA_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3777_elements(45) & convTransposeA_CP_3777_elements(47) & convTransposeA_CP_3777_elements(49);
      gj_convTransposeA_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3777_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	68 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1734_final_index_sum_regn_sample_complete
      -- CP-element group 59: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1734_final_index_sum_regn_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1734_final_index_sum_regn_Sample/ack
      -- 
    ack_4281_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1734_index_offset_ack_0, ack => convTransposeA_CP_3777_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	102 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (11) 
      -- CP-element group 60: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/addr_of_1735_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1734_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1734_offset_calculated
      -- CP-element group 60: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1734_final_index_sum_regn_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1734_final_index_sum_regn_Update/ack
      -- CP-element group 60: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1734_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1734_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1734_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1734_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/addr_of_1735_request/$entry
      -- CP-element group 60: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/addr_of_1735_request/req
      -- 
    ack_4286_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1734_index_offset_ack_1, ack => convTransposeA_CP_3777_elements(60)); -- 
    req_4295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(60), ack => addr_of_1735_final_reg_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/addr_of_1735_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/addr_of_1735_request/$exit
      -- CP-element group 61: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/addr_of_1735_request/ack
      -- 
    ack_4296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1735_final_reg_ack_0, ack => convTransposeA_CP_3777_elements(61)); -- 
    -- CP-element group 62:  fork  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	102 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (19) 
      -- CP-element group 62: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/addr_of_1735_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/addr_of_1735_complete/$exit
      -- CP-element group 62: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/addr_of_1735_complete/ack
      -- CP-element group 62: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1738_base_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1738_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1738_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1738_base_address_resized
      -- CP-element group 62: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1738_base_addr_resize/$entry
      -- CP-element group 62: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1738_base_addr_resize/$exit
      -- CP-element group 62: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1738_base_addr_resize/base_resize_req
      -- CP-element group 62: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1738_base_addr_resize/base_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1738_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1738_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1738_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1738_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1738_word_addrgen/$entry
      -- CP-element group 62: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1738_word_addrgen/$exit
      -- CP-element group 62: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1738_word_addrgen/root_register_req
      -- CP-element group 62: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1738_word_addrgen/root_register_ack
      -- 
    ack_4301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1735_final_reg_ack_1, ack => convTransposeA_CP_3777_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1738_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1738_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1738_Sample/ptr_deref_1738_Split/$entry
      -- CP-element group 63: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1738_Sample/ptr_deref_1738_Split/$exit
      -- CP-element group 63: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1738_Sample/ptr_deref_1738_Split/split_req
      -- CP-element group 63: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1738_Sample/ptr_deref_1738_Split/split_ack
      -- CP-element group 63: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1738_Sample/word_access_start/$entry
      -- CP-element group 63: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1738_Sample/word_access_start/word_0/$entry
      -- CP-element group 63: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1738_Sample/word_access_start/word_0/rr
      -- 
    rr_4339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(63), ack => ptr_deref_1738_store_0_req_0); -- 
    convTransposeA_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3777_elements(57) & convTransposeA_CP_3777_elements(62);
      gj_convTransposeA_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3777_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1738_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1738_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1738_Sample/word_access_start/$exit
      -- CP-element group 64: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1738_Sample/word_access_start/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1738_Sample/word_access_start/word_0/ra
      -- 
    ra_4340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1738_store_0_ack_0, ack => convTransposeA_CP_3777_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	102 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	68 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1738_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1738_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1738_Update/word_access_complete/$exit
      -- CP-element group 65: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1738_Update/word_access_complete/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1738_Update/word_access_complete/word_0/ca
      -- 
    ca_4351_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1738_store_0_ack_1, ack => convTransposeA_CP_3777_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	102 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1743_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1743_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1743_Sample/ra
      -- 
    ra_4360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1743_inst_ack_0, ack => convTransposeA_CP_3777_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	102 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1743_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1743_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1743_Update/ca
      -- 
    ca_4365_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1743_inst_ack_1, ack => convTransposeA_CP_3777_elements(67)); -- 
    -- CP-element group 68:  branch  join  transition  place  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	52 
    -- CP-element group 68: 	59 
    -- CP-element group 68: 	65 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (10) 
      -- CP-element group 68: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755__exit__
      -- CP-element group 68: 	 branch_block_stmt_1496/if_stmt_1756__entry__
      -- CP-element group 68: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/$exit
      -- CP-element group 68: 	 branch_block_stmt_1496/if_stmt_1756_dead_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1496/if_stmt_1756_eval_test/$entry
      -- CP-element group 68: 	 branch_block_stmt_1496/if_stmt_1756_eval_test/$exit
      -- CP-element group 68: 	 branch_block_stmt_1496/if_stmt_1756_eval_test/branch_req
      -- CP-element group 68: 	 branch_block_stmt_1496/R_cmp_1757_place
      -- CP-element group 68: 	 branch_block_stmt_1496/if_stmt_1756_if_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1496/if_stmt_1756_else_link/$entry
      -- 
    branch_req_4373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(68), ack => if_stmt_1756_branch_req_0); -- 
    convTransposeA_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3777_elements(52) & convTransposeA_CP_3777_elements(59) & convTransposeA_CP_3777_elements(65) & convTransposeA_CP_3777_elements(67);
      gj_convTransposeA_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3777_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	111 
    -- CP-element group 69: 	112 
    -- CP-element group 69: 	114 
    -- CP-element group 69: 	115 
    -- CP-element group 69: 	117 
    -- CP-element group 69: 	118 
    -- CP-element group 69:  members (40) 
      -- CP-element group 69: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1832/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1832/$entry
      -- CP-element group 69: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1814/phi_stmt_1814_sources/type_cast_1820/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1814/$entry
      -- CP-element group 69: 	 branch_block_stmt_1496/merge_stmt_1762__exit__
      -- CP-element group 69: 	 branch_block_stmt_1496/assign_stmt_1768__entry__
      -- CP-element group 69: 	 branch_block_stmt_1496/assign_stmt_1768__exit__
      -- CP-element group 69: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123
      -- CP-element group 69: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1832/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1814/phi_stmt_1814_sources/type_cast_1820/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1814/phi_stmt_1814_sources/type_cast_1820/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1496/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1814/phi_stmt_1814_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1496/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 69: 	 branch_block_stmt_1496/merge_stmt_1762_PhiAck/$entry
      -- CP-element group 69: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1832/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1827/$entry
      -- CP-element group 69: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1821/phi_stmt_1821_sources/type_cast_1824/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1821/phi_stmt_1821_sources/type_cast_1824/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1832/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1814/phi_stmt_1814_sources/type_cast_1820/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1821/phi_stmt_1821_sources/type_cast_1824/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1821/phi_stmt_1821_sources/type_cast_1824/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1821/phi_stmt_1821_sources/type_cast_1824/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1496/merge_stmt_1762_PhiReqMerge
      -- CP-element group 69: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1821/phi_stmt_1821_sources/type_cast_1824/$entry
      -- CP-element group 69: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1821/phi_stmt_1821_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1814/phi_stmt_1814_sources/type_cast_1820/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1832/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1814/phi_stmt_1814_sources/type_cast_1820/$entry
      -- CP-element group 69: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1821/$entry
      -- CP-element group 69: 	 branch_block_stmt_1496/merge_stmt_1762_PhiAck/dummy
      -- CP-element group 69: 	 branch_block_stmt_1496/merge_stmt_1762_PhiAck/$exit
      -- CP-element group 69: 	 branch_block_stmt_1496/if_stmt_1756_if_link/$exit
      -- CP-element group 69: 	 branch_block_stmt_1496/if_stmt_1756_if_link/if_choice_transition
      -- CP-element group 69: 	 branch_block_stmt_1496/whilex_xbody_ifx_xthen
      -- CP-element group 69: 	 branch_block_stmt_1496/assign_stmt_1768/$entry
      -- CP-element group 69: 	 branch_block_stmt_1496/assign_stmt_1768/$exit
      -- 
    if_choice_transition_4378_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1756_branch_ack_1, ack => convTransposeA_CP_3777_elements(69)); -- 
    cr_4700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(69), ack => type_cast_1832_inst_req_1); -- 
    rr_4741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(69), ack => type_cast_1820_inst_req_0); -- 
    cr_4746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(69), ack => type_cast_1820_inst_req_1); -- 
    cr_4723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(69), ack => type_cast_1824_inst_req_1); -- 
    rr_4718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(69), ack => type_cast_1824_inst_req_0); -- 
    rr_4695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(69), ack => type_cast_1832_inst_req_0); -- 
    -- CP-element group 70:  fork  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70: 	74 
    -- CP-element group 70:  members (21) 
      -- CP-element group 70: 	 branch_block_stmt_1496/merge_stmt_1770__exit__
      -- CP-element group 70: 	 branch_block_stmt_1496/assign_stmt_1776_to_assign_stmt_1806__entry__
      -- CP-element group 70: 	 branch_block_stmt_1496/merge_stmt_1770_PhiReqMerge
      -- CP-element group 70: 	 branch_block_stmt_1496/merge_stmt_1770_PhiAck/dummy
      -- CP-element group 70: 	 branch_block_stmt_1496/merge_stmt_1770_PhiAck/$exit
      -- CP-element group 70: 	 branch_block_stmt_1496/merge_stmt_1770_PhiAck/$entry
      -- CP-element group 70: 	 branch_block_stmt_1496/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 70: 	 branch_block_stmt_1496/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_1496/if_stmt_1756_else_link/$exit
      -- CP-element group 70: 	 branch_block_stmt_1496/if_stmt_1756_else_link/else_choice_transition
      -- CP-element group 70: 	 branch_block_stmt_1496/whilex_xbody_ifx_xelse
      -- CP-element group 70: 	 branch_block_stmt_1496/assign_stmt_1776_to_assign_stmt_1806/$entry
      -- CP-element group 70: 	 branch_block_stmt_1496/assign_stmt_1776_to_assign_stmt_1806/type_cast_1784_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_1496/assign_stmt_1776_to_assign_stmt_1806/type_cast_1784_update_start_
      -- CP-element group 70: 	 branch_block_stmt_1496/assign_stmt_1776_to_assign_stmt_1806/type_cast_1784_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_1496/assign_stmt_1776_to_assign_stmt_1806/type_cast_1784_Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_1496/assign_stmt_1776_to_assign_stmt_1806/type_cast_1784_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1496/assign_stmt_1776_to_assign_stmt_1806/type_cast_1784_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_1496/assign_stmt_1776_to_assign_stmt_1806/type_cast_1800_update_start_
      -- CP-element group 70: 	 branch_block_stmt_1496/assign_stmt_1776_to_assign_stmt_1806/type_cast_1800_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1496/assign_stmt_1776_to_assign_stmt_1806/type_cast_1800_Update/cr
      -- 
    else_choice_transition_4382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1756_branch_ack_0, ack => convTransposeA_CP_3777_elements(70)); -- 
    rr_4398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(70), ack => type_cast_1784_inst_req_0); -- 
    cr_4403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(70), ack => type_cast_1784_inst_req_1); -- 
    cr_4417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(70), ack => type_cast_1800_inst_req_1); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_1496/assign_stmt_1776_to_assign_stmt_1806/type_cast_1784_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_1496/assign_stmt_1776_to_assign_stmt_1806/type_cast_1784_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_1496/assign_stmt_1776_to_assign_stmt_1806/type_cast_1784_Sample/ra
      -- 
    ra_4399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1784_inst_ack_0, ack => convTransposeA_CP_3777_elements(71)); -- 
    -- CP-element group 72:  transition  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (6) 
      -- CP-element group 72: 	 branch_block_stmt_1496/assign_stmt_1776_to_assign_stmt_1806/type_cast_1784_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_1496/assign_stmt_1776_to_assign_stmt_1806/type_cast_1784_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_1496/assign_stmt_1776_to_assign_stmt_1806/type_cast_1784_Update/ca
      -- CP-element group 72: 	 branch_block_stmt_1496/assign_stmt_1776_to_assign_stmt_1806/type_cast_1800_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_1496/assign_stmt_1776_to_assign_stmt_1806/type_cast_1800_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_1496/assign_stmt_1776_to_assign_stmt_1806/type_cast_1800_Sample/rr
      -- 
    ca_4404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1784_inst_ack_1, ack => convTransposeA_CP_3777_elements(72)); -- 
    rr_4412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(72), ack => type_cast_1800_inst_req_0); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1496/assign_stmt_1776_to_assign_stmt_1806/type_cast_1800_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_1496/assign_stmt_1776_to_assign_stmt_1806/type_cast_1800_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_1496/assign_stmt_1776_to_assign_stmt_1806/type_cast_1800_Sample/ra
      -- 
    ra_4413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1800_inst_ack_0, ack => convTransposeA_CP_3777_elements(73)); -- 
    -- CP-element group 74:  branch  transition  place  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	70 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (13) 
      -- CP-element group 74: 	 branch_block_stmt_1496/assign_stmt_1776_to_assign_stmt_1806__exit__
      -- CP-element group 74: 	 branch_block_stmt_1496/if_stmt_1807__entry__
      -- CP-element group 74: 	 branch_block_stmt_1496/assign_stmt_1776_to_assign_stmt_1806/$exit
      -- CP-element group 74: 	 branch_block_stmt_1496/assign_stmt_1776_to_assign_stmt_1806/type_cast_1800_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_1496/assign_stmt_1776_to_assign_stmt_1806/type_cast_1800_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_1496/assign_stmt_1776_to_assign_stmt_1806/type_cast_1800_Update/ca
      -- CP-element group 74: 	 branch_block_stmt_1496/if_stmt_1807_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1496/if_stmt_1807_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_1496/if_stmt_1807_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_1496/if_stmt_1807_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_1496/R_cmp112_1808_place
      -- CP-element group 74: 	 branch_block_stmt_1496/if_stmt_1807_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1496/if_stmt_1807_else_link/$entry
      -- 
    ca_4418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1800_inst_ack_1, ack => convTransposeA_CP_3777_elements(74)); -- 
    branch_req_4426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(74), ack => if_stmt_1807_branch_req_0); -- 
    -- CP-element group 75:  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (15) 
      -- CP-element group 75: 	 branch_block_stmt_1496/merge_stmt_1841__exit__
      -- CP-element group 75: 	 branch_block_stmt_1496/assign_stmt_1846__entry__
      -- CP-element group 75: 	 branch_block_stmt_1496/merge_stmt_1841_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_1496/merge_stmt_1841_PhiAck/dummy
      -- CP-element group 75: 	 branch_block_stmt_1496/merge_stmt_1841_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_1496/merge_stmt_1841_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_1496/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_1496/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_1496/assign_stmt_1846/WPIPE_Block0_done_1843_Sample/req
      -- CP-element group 75: 	 branch_block_stmt_1496/assign_stmt_1846/WPIPE_Block0_done_1843_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_1496/if_stmt_1807_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_1496/if_stmt_1807_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_1496/ifx_xelse_whilex_xend
      -- CP-element group 75: 	 branch_block_stmt_1496/assign_stmt_1846/$entry
      -- CP-element group 75: 	 branch_block_stmt_1496/assign_stmt_1846/WPIPE_Block0_done_1843_sample_start_
      -- 
    if_choice_transition_4431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1807_branch_ack_1, ack => convTransposeA_CP_3777_elements(75)); -- 
    req_4451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(75), ack => WPIPE_Block0_done_1843_inst_req_0); -- 
    -- CP-element group 76:  fork  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	103 
    -- CP-element group 76: 	104 
    -- CP-element group 76: 	106 
    -- CP-element group 76: 	107 
    -- CP-element group 76: 	109 
    -- CP-element group 76:  members (22) 
      -- CP-element group 76: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1821/$entry
      -- CP-element group 76: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1830/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1830/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1830/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1830/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1814/phi_stmt_1814_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1830/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1814/$entry
      -- CP-element group 76: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1830/$entry
      -- CP-element group 76: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1821/phi_stmt_1821_sources/type_cast_1826/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1821/phi_stmt_1821_sources/type_cast_1826/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1827/$entry
      -- CP-element group 76: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1821/phi_stmt_1821_sources/type_cast_1826/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1821/phi_stmt_1821_sources/type_cast_1826/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1821/phi_stmt_1821_sources/type_cast_1826/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1821/phi_stmt_1821_sources/type_cast_1826/$entry
      -- CP-element group 76: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1821/phi_stmt_1821_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1496/if_stmt_1807_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_1496/if_stmt_1807_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123
      -- 
    else_choice_transition_4435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1807_branch_ack_0, ack => convTransposeA_CP_3777_elements(76)); -- 
    cr_4643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(76), ack => type_cast_1830_inst_req_1); -- 
    rr_4638_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4638_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(76), ack => type_cast_1830_inst_req_0); -- 
    cr_4666_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4666_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(76), ack => type_cast_1826_inst_req_1); -- 
    rr_4661_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4661_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(76), ack => type_cast_1826_inst_req_0); -- 
    -- CP-element group 77:  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (6) 
      -- CP-element group 77: 	 branch_block_stmt_1496/assign_stmt_1846/WPIPE_Block0_done_1843_Update/req
      -- CP-element group 77: 	 branch_block_stmt_1496/assign_stmt_1846/WPIPE_Block0_done_1843_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_1496/assign_stmt_1846/WPIPE_Block0_done_1843_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1496/assign_stmt_1846/WPIPE_Block0_done_1843_Sample/ack
      -- CP-element group 77: 	 branch_block_stmt_1496/assign_stmt_1846/WPIPE_Block0_done_1843_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_1496/assign_stmt_1846/WPIPE_Block0_done_1843_update_start_
      -- 
    ack_4452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1843_inst_ack_0, ack => convTransposeA_CP_3777_elements(77)); -- 
    req_4456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(77), ack => WPIPE_Block0_done_1843_inst_req_1); -- 
    -- CP-element group 78:  transition  place  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (16) 
      -- CP-element group 78: 	 branch_block_stmt_1496/$exit
      -- CP-element group 78: 	 branch_block_stmt_1496/merge_stmt_1848__exit__
      -- CP-element group 78: 	 branch_block_stmt_1496/assign_stmt_1846__exit__
      -- CP-element group 78: 	 branch_block_stmt_1496/assign_stmt_1846/WPIPE_Block0_done_1843_Update/ack
      -- CP-element group 78: 	 branch_block_stmt_1496/branch_block_stmt_1496__exit__
      -- CP-element group 78: 	 branch_block_stmt_1496/return__
      -- CP-element group 78: 	 $exit
      -- CP-element group 78: 	 branch_block_stmt_1496/merge_stmt_1848_PhiReqMerge
      -- CP-element group 78: 	 branch_block_stmt_1496/merge_stmt_1848_PhiAck/dummy
      -- CP-element group 78: 	 branch_block_stmt_1496/merge_stmt_1848_PhiAck/$exit
      -- CP-element group 78: 	 branch_block_stmt_1496/merge_stmt_1848_PhiAck/$entry
      -- CP-element group 78: 	 branch_block_stmt_1496/return___PhiReq/$exit
      -- CP-element group 78: 	 branch_block_stmt_1496/return___PhiReq/$entry
      -- CP-element group 78: 	 branch_block_stmt_1496/assign_stmt_1846/WPIPE_Block0_done_1843_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_1496/assign_stmt_1846/$exit
      -- CP-element group 78: 	 branch_block_stmt_1496/assign_stmt_1846/WPIPE_Block0_done_1843_update_completed_
      -- 
    ack_4457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1843_inst_ack_1, ack => convTransposeA_CP_3777_elements(78)); -- 
    -- CP-element group 79:  transition  output  delay-element  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	43 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	83 
    -- CP-element group 79:  members (4) 
      -- CP-element group 79: 	 branch_block_stmt_1496/entry_whilex_xbody_PhiReq/phi_stmt_1605/$exit
      -- CP-element group 79: 	 branch_block_stmt_1496/entry_whilex_xbody_PhiReq/phi_stmt_1605/phi_stmt_1605_sources/$exit
      -- CP-element group 79: 	 branch_block_stmt_1496/entry_whilex_xbody_PhiReq/phi_stmt_1605/phi_stmt_1605_sources/type_cast_1609_konst_delay_trans
      -- CP-element group 79: 	 branch_block_stmt_1496/entry_whilex_xbody_PhiReq/phi_stmt_1605/phi_stmt_1605_req
      -- 
    phi_stmt_1605_req_4468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1605_req_4468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(79), ack => phi_stmt_1605_req_0); -- 
    -- Element group convTransposeA_CP_3777_elements(79) is a control-delay.
    cp_element_79_delay: control_delay_element  generic map(name => " 79_delay", delay_value => 1)  port map(req => convTransposeA_CP_3777_elements(43), ack => convTransposeA_CP_3777_elements(79), clk => clk, reset =>reset);
    -- CP-element group 80:  transition  output  delay-element  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	43 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	83 
    -- CP-element group 80:  members (4) 
      -- CP-element group 80: 	 branch_block_stmt_1496/entry_whilex_xbody_PhiReq/phi_stmt_1612/phi_stmt_1612_sources/$exit
      -- CP-element group 80: 	 branch_block_stmt_1496/entry_whilex_xbody_PhiReq/phi_stmt_1612/phi_stmt_1612_sources/type_cast_1616_konst_delay_trans
      -- CP-element group 80: 	 branch_block_stmt_1496/entry_whilex_xbody_PhiReq/phi_stmt_1612/phi_stmt_1612_req
      -- CP-element group 80: 	 branch_block_stmt_1496/entry_whilex_xbody_PhiReq/phi_stmt_1612/$exit
      -- 
    phi_stmt_1612_req_4476_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1612_req_4476_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(80), ack => phi_stmt_1612_req_0); -- 
    -- Element group convTransposeA_CP_3777_elements(80) is a control-delay.
    cp_element_80_delay: control_delay_element  generic map(name => " 80_delay", delay_value => 1)  port map(req => convTransposeA_CP_3777_elements(43), ack => convTransposeA_CP_3777_elements(80), clk => clk, reset =>reset);
    -- CP-element group 81:  transition  output  delay-element  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	43 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (4) 
      -- CP-element group 81: 	 branch_block_stmt_1496/entry_whilex_xbody_PhiReq/phi_stmt_1619/phi_stmt_1619_req
      -- CP-element group 81: 	 branch_block_stmt_1496/entry_whilex_xbody_PhiReq/phi_stmt_1619/phi_stmt_1619_sources/type_cast_1623_konst_delay_trans
      -- CP-element group 81: 	 branch_block_stmt_1496/entry_whilex_xbody_PhiReq/phi_stmt_1619/phi_stmt_1619_sources/$exit
      -- CP-element group 81: 	 branch_block_stmt_1496/entry_whilex_xbody_PhiReq/phi_stmt_1619/$exit
      -- 
    phi_stmt_1619_req_4484_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1619_req_4484_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(81), ack => phi_stmt_1619_req_0); -- 
    -- Element group convTransposeA_CP_3777_elements(81) is a control-delay.
    cp_element_81_delay: control_delay_element  generic map(name => " 81_delay", delay_value => 1)  port map(req => convTransposeA_CP_3777_elements(43), ack => convTransposeA_CP_3777_elements(81), clk => clk, reset =>reset);
    -- CP-element group 82:  transition  output  delay-element  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	43 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (4) 
      -- CP-element group 82: 	 branch_block_stmt_1496/entry_whilex_xbody_PhiReq/phi_stmt_1626/phi_stmt_1626_sources/type_cast_1630_konst_delay_trans
      -- CP-element group 82: 	 branch_block_stmt_1496/entry_whilex_xbody_PhiReq/phi_stmt_1626/phi_stmt_1626_sources/$exit
      -- CP-element group 82: 	 branch_block_stmt_1496/entry_whilex_xbody_PhiReq/phi_stmt_1626/phi_stmt_1626_req
      -- CP-element group 82: 	 branch_block_stmt_1496/entry_whilex_xbody_PhiReq/phi_stmt_1626/$exit
      -- 
    phi_stmt_1626_req_4492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1626_req_4492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(82), ack => phi_stmt_1626_req_0); -- 
    -- Element group convTransposeA_CP_3777_elements(82) is a control-delay.
    cp_element_82_delay: control_delay_element  generic map(name => " 82_delay", delay_value => 1)  port map(req => convTransposeA_CP_3777_elements(43), ack => convTransposeA_CP_3777_elements(82), clk => clk, reset =>reset);
    -- CP-element group 83:  join  transition  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	79 
    -- CP-element group 83: 	80 
    -- CP-element group 83: 	81 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	97 
    -- CP-element group 83:  members (1) 
      -- CP-element group 83: 	 branch_block_stmt_1496/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3777_elements(79) & convTransposeA_CP_3777_elements(80) & convTransposeA_CP_3777_elements(81) & convTransposeA_CP_3777_elements(82);
      gj_convTransposeA_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3777_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	1 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1605/phi_stmt_1605_sources/type_cast_1611/SplitProtocol/Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1605/phi_stmt_1605_sources/type_cast_1611/SplitProtocol/Sample/ra
      -- 
    ra_4512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1611_inst_ack_0, ack => convTransposeA_CP_3777_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	1 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1605/phi_stmt_1605_sources/type_cast_1611/SplitProtocol/Update/ca
      -- CP-element group 85: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1605/phi_stmt_1605_sources/type_cast_1611/SplitProtocol/Update/$exit
      -- 
    ca_4517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1611_inst_ack_1, ack => convTransposeA_CP_3777_elements(85)); -- 
    -- CP-element group 86:  join  transition  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	96 
    -- CP-element group 86:  members (5) 
      -- CP-element group 86: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1605/$exit
      -- CP-element group 86: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1605/phi_stmt_1605_sources/$exit
      -- CP-element group 86: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1605/phi_stmt_1605_sources/type_cast_1611/$exit
      -- CP-element group 86: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1605/phi_stmt_1605_sources/type_cast_1611/SplitProtocol/$exit
      -- CP-element group 86: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1605/phi_stmt_1605_req
      -- 
    phi_stmt_1605_req_4518_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1605_req_4518_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(86), ack => phi_stmt_1605_req_1); -- 
    convTransposeA_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3777_elements(84) & convTransposeA_CP_3777_elements(85);
      gj_convTransposeA_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3777_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	1 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1612/phi_stmt_1612_sources/type_cast_1618/SplitProtocol/Sample/ra
      -- CP-element group 87: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1612/phi_stmt_1612_sources/type_cast_1618/SplitProtocol/Sample/$exit
      -- 
    ra_4535_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1618_inst_ack_0, ack => convTransposeA_CP_3777_elements(87)); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	1 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1612/phi_stmt_1612_sources/type_cast_1618/SplitProtocol/Update/ca
      -- CP-element group 88: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1612/phi_stmt_1612_sources/type_cast_1618/SplitProtocol/Update/$exit
      -- 
    ca_4540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1618_inst_ack_1, ack => convTransposeA_CP_3777_elements(88)); -- 
    -- CP-element group 89:  join  transition  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	96 
    -- CP-element group 89:  members (5) 
      -- CP-element group 89: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1612/phi_stmt_1612_req
      -- CP-element group 89: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1612/phi_stmt_1612_sources/type_cast_1618/SplitProtocol/$exit
      -- CP-element group 89: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1612/phi_stmt_1612_sources/type_cast_1618/$exit
      -- CP-element group 89: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1612/phi_stmt_1612_sources/$exit
      -- CP-element group 89: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1612/$exit
      -- 
    phi_stmt_1612_req_4541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1612_req_4541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(89), ack => phi_stmt_1612_req_1); -- 
    convTransposeA_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3777_elements(87) & convTransposeA_CP_3777_elements(88);
      gj_convTransposeA_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3777_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	1 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1619/phi_stmt_1619_sources/type_cast_1625/SplitProtocol/Sample/ra
      -- CP-element group 90: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1619/phi_stmt_1619_sources/type_cast_1625/SplitProtocol/Sample/$exit
      -- 
    ra_4558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1625_inst_ack_0, ack => convTransposeA_CP_3777_elements(90)); -- 
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	1 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1619/phi_stmt_1619_sources/type_cast_1625/SplitProtocol/Update/ca
      -- CP-element group 91: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1619/phi_stmt_1619_sources/type_cast_1625/SplitProtocol/Update/$exit
      -- 
    ca_4563_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1625_inst_ack_1, ack => convTransposeA_CP_3777_elements(91)); -- 
    -- CP-element group 92:  join  transition  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	96 
    -- CP-element group 92:  members (5) 
      -- CP-element group 92: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1619/phi_stmt_1619_req
      -- CP-element group 92: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1619/phi_stmt_1619_sources/type_cast_1625/SplitProtocol/$exit
      -- CP-element group 92: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1619/phi_stmt_1619_sources/type_cast_1625/$exit
      -- CP-element group 92: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1619/phi_stmt_1619_sources/$exit
      -- CP-element group 92: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1619/$exit
      -- 
    phi_stmt_1619_req_4564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1619_req_4564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(92), ack => phi_stmt_1619_req_1); -- 
    convTransposeA_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3777_elements(90) & convTransposeA_CP_3777_elements(91);
      gj_convTransposeA_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3777_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	1 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1626/phi_stmt_1626_sources/type_cast_1632/SplitProtocol/Sample/ra
      -- CP-element group 93: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1626/phi_stmt_1626_sources/type_cast_1632/SplitProtocol/Sample/$exit
      -- 
    ra_4581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1632_inst_ack_0, ack => convTransposeA_CP_3777_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	1 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1626/phi_stmt_1626_sources/type_cast_1632/SplitProtocol/Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1626/phi_stmt_1626_sources/type_cast_1632/SplitProtocol/Update/ca
      -- 
    ca_4586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1632_inst_ack_1, ack => convTransposeA_CP_3777_elements(94)); -- 
    -- CP-element group 95:  join  transition  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (5) 
      -- CP-element group 95: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1626/phi_stmt_1626_sources/type_cast_1632/SplitProtocol/$exit
      -- CP-element group 95: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1626/phi_stmt_1626_sources/type_cast_1632/$exit
      -- CP-element group 95: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1626/phi_stmt_1626_sources/$exit
      -- CP-element group 95: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1626/$exit
      -- CP-element group 95: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1626/phi_stmt_1626_req
      -- 
    phi_stmt_1626_req_4587_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1626_req_4587_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(95), ack => phi_stmt_1626_req_1); -- 
    convTransposeA_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3777_elements(93) & convTransposeA_CP_3777_elements(94);
      gj_convTransposeA_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3777_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  join  transition  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	86 
    -- CP-element group 96: 	89 
    -- CP-element group 96: 	92 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_1496/ifx_xend123_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3777_elements(86) & convTransposeA_CP_3777_elements(89) & convTransposeA_CP_3777_elements(92) & convTransposeA_CP_3777_elements(95);
      gj_convTransposeA_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3777_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  merge  fork  transition  place  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	83 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97: 	99 
    -- CP-element group 97: 	100 
    -- CP-element group 97: 	101 
    -- CP-element group 97:  members (2) 
      -- CP-element group 97: 	 branch_block_stmt_1496/merge_stmt_1604_PhiAck/$entry
      -- CP-element group 97: 	 branch_block_stmt_1496/merge_stmt_1604_PhiReqMerge
      -- 
    convTransposeA_CP_3777_elements(97) <= OrReduce(convTransposeA_CP_3777_elements(83) & convTransposeA_CP_3777_elements(96));
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	102 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_1496/merge_stmt_1604_PhiAck/phi_stmt_1605_ack
      -- 
    phi_stmt_1605_ack_4592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1605_ack_0, ack => convTransposeA_CP_3777_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	97 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	102 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_1496/merge_stmt_1604_PhiAck/phi_stmt_1612_ack
      -- 
    phi_stmt_1612_ack_4593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1612_ack_0, ack => convTransposeA_CP_3777_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	97 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	102 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_1496/merge_stmt_1604_PhiAck/phi_stmt_1619_ack
      -- 
    phi_stmt_1619_ack_4594_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1619_ack_0, ack => convTransposeA_CP_3777_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	97 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	102 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_1496/merge_stmt_1604_PhiAck/phi_stmt_1626_ack
      -- 
    phi_stmt_1626_ack_4595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1626_ack_0, ack => convTransposeA_CP_3777_elements(101)); -- 
    -- CP-element group 102:  join  fork  transition  place  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	98 
    -- CP-element group 102: 	99 
    -- CP-element group 102: 	100 
    -- CP-element group 102: 	101 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	44 
    -- CP-element group 102: 	45 
    -- CP-element group 102: 	46 
    -- CP-element group 102: 	47 
    -- CP-element group 102: 	48 
    -- CP-element group 102: 	49 
    -- CP-element group 102: 	50 
    -- CP-element group 102: 	51 
    -- CP-element group 102: 	53 
    -- CP-element group 102: 	55 
    -- CP-element group 102: 	57 
    -- CP-element group 102: 	60 
    -- CP-element group 102: 	62 
    -- CP-element group 102: 	65 
    -- CP-element group 102: 	66 
    -- CP-element group 102: 	67 
    -- CP-element group 102:  members (56) 
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755__entry__
      -- CP-element group 102: 	 branch_block_stmt_1496/merge_stmt_1604__exit__
      -- CP-element group 102: 	 branch_block_stmt_1496/merge_stmt_1604_PhiAck/$exit
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/$entry
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1667_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1667_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1667_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1667_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1667_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1667_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1671_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1671_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1671_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1671_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1671_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1671_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1675_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1675_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1675_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1675_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1675_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1675_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1705_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1705_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1705_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1705_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1705_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1705_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/addr_of_1712_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1711_final_index_sum_regn_update_start
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1711_final_index_sum_regn_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1711_final_index_sum_regn_Update/req
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/addr_of_1712_complete/$entry
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/addr_of_1712_complete/req
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1716_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1716_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1716_Update/word_access_complete/$entry
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1716_Update/word_access_complete/word_0/$entry
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1716_Update/word_access_complete/word_0/cr
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/addr_of_1735_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1734_final_index_sum_regn_update_start
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1734_final_index_sum_regn_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/array_obj_ref_1734_final_index_sum_regn_Update/req
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/addr_of_1735_complete/$entry
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/addr_of_1735_complete/req
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1738_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1738_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1738_Update/word_access_complete/$entry
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1738_Update/word_access_complete/word_0/$entry
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/ptr_deref_1738_Update/word_access_complete/word_0/cr
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1743_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1743_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1743_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1743_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1743_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1496/assign_stmt_1639_to_assign_stmt_1755/type_cast_1743_Update/cr
      -- 
    rr_4111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(102), ack => type_cast_1667_inst_req_0); -- 
    cr_4116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(102), ack => type_cast_1667_inst_req_1); -- 
    rr_4125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(102), ack => type_cast_1671_inst_req_0); -- 
    cr_4130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(102), ack => type_cast_1671_inst_req_1); -- 
    rr_4139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(102), ack => type_cast_1675_inst_req_0); -- 
    cr_4144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(102), ack => type_cast_1675_inst_req_1); -- 
    rr_4153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(102), ack => type_cast_1705_inst_req_0); -- 
    cr_4158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(102), ack => type_cast_1705_inst_req_1); -- 
    req_4189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(102), ack => array_obj_ref_1711_index_offset_req_1); -- 
    req_4204_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4204_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(102), ack => addr_of_1712_final_reg_req_1); -- 
    cr_4249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(102), ack => ptr_deref_1716_load_0_req_1); -- 
    req_4285_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4285_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(102), ack => array_obj_ref_1734_index_offset_req_1); -- 
    req_4300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(102), ack => addr_of_1735_final_reg_req_1); -- 
    cr_4350_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4350_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(102), ack => ptr_deref_1738_store_0_req_1); -- 
    rr_4359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(102), ack => type_cast_1743_inst_req_0); -- 
    cr_4364_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4364_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(102), ack => type_cast_1743_inst_req_1); -- 
    convTransposeA_cp_element_group_102: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_102"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3777_elements(98) & convTransposeA_CP_3777_elements(99) & convTransposeA_CP_3777_elements(100) & convTransposeA_CP_3777_elements(101);
      gj_convTransposeA_cp_element_group_102 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3777_elements(102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	76 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	105 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1830/SplitProtocol/Sample/ra
      -- CP-element group 103: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1830/SplitProtocol/Sample/$exit
      -- 
    ra_4639_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1830_inst_ack_0, ack => convTransposeA_CP_3777_elements(103)); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	76 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1830/SplitProtocol/Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1830/SplitProtocol/Update/ca
      -- 
    ca_4644_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1830_inst_ack_1, ack => convTransposeA_CP_3777_elements(104)); -- 
    -- CP-element group 105:  join  transition  output  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	103 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	110 
    -- CP-element group 105:  members (5) 
      -- CP-element group 105: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_req
      -- CP-element group 105: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1830/SplitProtocol/$exit
      -- CP-element group 105: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1830/$exit
      -- CP-element group 105: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/$exit
      -- CP-element group 105: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1827/$exit
      -- 
    phi_stmt_1827_req_4645_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1827_req_4645_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(105), ack => phi_stmt_1827_req_0); -- 
    convTransposeA_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3777_elements(103) & convTransposeA_CP_3777_elements(104);
      gj_convTransposeA_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3777_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	76 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1821/phi_stmt_1821_sources/type_cast_1826/SplitProtocol/Sample/ra
      -- CP-element group 106: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1821/phi_stmt_1821_sources/type_cast_1826/SplitProtocol/Sample/$exit
      -- 
    ra_4662_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1826_inst_ack_0, ack => convTransposeA_CP_3777_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	76 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1821/phi_stmt_1821_sources/type_cast_1826/SplitProtocol/Update/ca
      -- CP-element group 107: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1821/phi_stmt_1821_sources/type_cast_1826/SplitProtocol/Update/$exit
      -- 
    ca_4667_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1826_inst_ack_1, ack => convTransposeA_CP_3777_elements(107)); -- 
    -- CP-element group 108:  join  transition  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	110 
    -- CP-element group 108:  members (5) 
      -- CP-element group 108: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1821/$exit
      -- CP-element group 108: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1821/phi_stmt_1821_req
      -- CP-element group 108: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1821/phi_stmt_1821_sources/type_cast_1826/SplitProtocol/$exit
      -- CP-element group 108: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1821/phi_stmt_1821_sources/type_cast_1826/$exit
      -- CP-element group 108: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1821/phi_stmt_1821_sources/$exit
      -- 
    phi_stmt_1821_req_4668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1821_req_4668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(108), ack => phi_stmt_1821_req_1); -- 
    convTransposeA_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3777_elements(106) & convTransposeA_CP_3777_elements(107);
      gj_convTransposeA_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3777_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  transition  output  delay-element  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	76 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109:  members (4) 
      -- CP-element group 109: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1814/phi_stmt_1814_req
      -- CP-element group 109: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1814/phi_stmt_1814_sources/type_cast_1818_konst_delay_trans
      -- CP-element group 109: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1814/phi_stmt_1814_sources/$exit
      -- CP-element group 109: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1814/$exit
      -- 
    phi_stmt_1814_req_4676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1814_req_4676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(109), ack => phi_stmt_1814_req_0); -- 
    -- Element group convTransposeA_CP_3777_elements(109) is a control-delay.
    cp_element_109_delay: control_delay_element  generic map(name => " 109_delay", delay_value => 1)  port map(req => convTransposeA_CP_3777_elements(76), ack => convTransposeA_CP_3777_elements(109), clk => clk, reset =>reset);
    -- CP-element group 110:  join  transition  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	105 
    -- CP-element group 110: 	108 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	121 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_1496/ifx_xelse_ifx_xend123_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3777_elements(105) & convTransposeA_CP_3777_elements(108) & convTransposeA_CP_3777_elements(109);
      gj_convTransposeA_cp_element_group_110 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3777_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	69 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	113 
    -- CP-element group 111:  members (2) 
      -- CP-element group 111: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1832/SplitProtocol/Sample/ra
      -- CP-element group 111: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1832/SplitProtocol/Sample/$exit
      -- 
    ra_4696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1832_inst_ack_0, ack => convTransposeA_CP_3777_elements(111)); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	69 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (2) 
      -- CP-element group 112: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1832/SplitProtocol/Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1832/SplitProtocol/Update/ca
      -- 
    ca_4701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1832_inst_ack_1, ack => convTransposeA_CP_3777_elements(112)); -- 
    -- CP-element group 113:  join  transition  output  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	111 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	120 
    -- CP-element group 113:  members (5) 
      -- CP-element group 113: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1832/$exit
      -- CP-element group 113: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1832/SplitProtocol/$exit
      -- CP-element group 113: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1827/$exit
      -- CP-element group 113: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/$exit
      -- CP-element group 113: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_req
      -- 
    phi_stmt_1827_req_4702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1827_req_4702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(113), ack => phi_stmt_1827_req_1); -- 
    convTransposeA_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3777_elements(111) & convTransposeA_CP_3777_elements(112);
      gj_convTransposeA_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3777_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	69 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (2) 
      -- CP-element group 114: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1821/phi_stmt_1821_sources/type_cast_1824/SplitProtocol/Sample/ra
      -- CP-element group 114: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1821/phi_stmt_1821_sources/type_cast_1824/SplitProtocol/Sample/$exit
      -- 
    ra_4719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1824_inst_ack_0, ack => convTransposeA_CP_3777_elements(114)); -- 
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	69 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1821/phi_stmt_1821_sources/type_cast_1824/SplitProtocol/Update/ca
      -- CP-element group 115: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1821/phi_stmt_1821_sources/type_cast_1824/SplitProtocol/Update/$exit
      -- 
    ca_4724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1824_inst_ack_1, ack => convTransposeA_CP_3777_elements(115)); -- 
    -- CP-element group 116:  join  transition  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	120 
    -- CP-element group 116:  members (5) 
      -- CP-element group 116: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1821/phi_stmt_1821_req
      -- CP-element group 116: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1821/phi_stmt_1821_sources/type_cast_1824/SplitProtocol/$exit
      -- CP-element group 116: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1821/phi_stmt_1821_sources/type_cast_1824/$exit
      -- CP-element group 116: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1821/phi_stmt_1821_sources/$exit
      -- CP-element group 116: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1821/$exit
      -- 
    phi_stmt_1821_req_4725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1821_req_4725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(116), ack => phi_stmt_1821_req_0); -- 
    convTransposeA_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3777_elements(114) & convTransposeA_CP_3777_elements(115);
      gj_convTransposeA_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3777_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	69 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	119 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1814/phi_stmt_1814_sources/type_cast_1820/SplitProtocol/Sample/ra
      -- CP-element group 117: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1814/phi_stmt_1814_sources/type_cast_1820/SplitProtocol/Sample/$exit
      -- 
    ra_4742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1820_inst_ack_0, ack => convTransposeA_CP_3777_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	69 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (2) 
      -- CP-element group 118: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1814/phi_stmt_1814_sources/type_cast_1820/SplitProtocol/Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1814/phi_stmt_1814_sources/type_cast_1820/SplitProtocol/Update/ca
      -- 
    ca_4747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1820_inst_ack_1, ack => convTransposeA_CP_3777_elements(118)); -- 
    -- CP-element group 119:  join  transition  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	117 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (5) 
      -- CP-element group 119: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1814/$exit
      -- CP-element group 119: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1814/phi_stmt_1814_req
      -- CP-element group 119: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1814/phi_stmt_1814_sources/type_cast_1820/SplitProtocol/$exit
      -- CP-element group 119: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1814/phi_stmt_1814_sources/type_cast_1820/$exit
      -- CP-element group 119: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1814/phi_stmt_1814_sources/$exit
      -- 
    phi_stmt_1814_req_4748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1814_req_4748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(119), ack => phi_stmt_1814_req_1); -- 
    convTransposeA_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3777_elements(117) & convTransposeA_CP_3777_elements(118);
      gj_convTransposeA_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3777_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  join  transition  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	113 
    -- CP-element group 120: 	116 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_1496/ifx_xthen_ifx_xend123_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3777_elements(113) & convTransposeA_CP_3777_elements(116) & convTransposeA_CP_3777_elements(119);
      gj_convTransposeA_cp_element_group_120 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3777_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  merge  fork  transition  place  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	110 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121: 	123 
    -- CP-element group 121: 	124 
    -- CP-element group 121:  members (2) 
      -- CP-element group 121: 	 branch_block_stmt_1496/merge_stmt_1813_PhiAck/$entry
      -- CP-element group 121: 	 branch_block_stmt_1496/merge_stmt_1813_PhiReqMerge
      -- 
    convTransposeA_CP_3777_elements(121) <= OrReduce(convTransposeA_CP_3777_elements(110) & convTransposeA_CP_3777_elements(120));
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	125 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_1496/merge_stmt_1813_PhiAck/phi_stmt_1814_ack
      -- 
    phi_stmt_1814_ack_4753_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1814_ack_0, ack => convTransposeA_CP_3777_elements(122)); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	121 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	125 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_1496/merge_stmt_1813_PhiAck/phi_stmt_1821_ack
      -- 
    phi_stmt_1821_ack_4754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1821_ack_0, ack => convTransposeA_CP_3777_elements(123)); -- 
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	121 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	125 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_1496/merge_stmt_1813_PhiAck/phi_stmt_1827_ack
      -- 
    phi_stmt_1827_ack_4755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1827_ack_0, ack => convTransposeA_CP_3777_elements(124)); -- 
    -- CP-element group 125:  join  transition  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	122 
    -- CP-element group 125: 	123 
    -- CP-element group 125: 	124 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	1 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_1496/merge_stmt_1813_PhiAck/$exit
      -- 
    convTransposeA_cp_element_group_125: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_125"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3777_elements(122) & convTransposeA_CP_3777_elements(123) & convTransposeA_CP_3777_elements(124);
      gj_convTransposeA_cp_element_group_125 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3777_elements(125), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom81_1733_resized : std_logic_vector(13 downto 0);
    signal R_idxprom81_1733_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_1710_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_1710_scaled : std_logic_vector(13 downto 0);
    signal add41_1564 : std_logic_vector(15 downto 0);
    signal add54_1575 : std_logic_vector(15 downto 0);
    signal add73_1686 : std_logic_vector(63 downto 0);
    signal add75_1696 : std_logic_vector(63 downto 0);
    signal add86_1750 : std_logic_vector(31 downto 0);
    signal add93_1768 : std_logic_vector(15 downto 0);
    signal add_1548 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_1644 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1711_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1711_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1711_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1711_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1711_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1711_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1734_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1734_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1734_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1734_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1734_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1734_root_address : std_logic_vector(13 downto 0);
    signal arrayidx77_1713 : std_logic_vector(31 downto 0);
    signal arrayidx82_1736 : std_logic_vector(31 downto 0);
    signal call11_1517 : std_logic_vector(15 downto 0);
    signal call13_1520 : std_logic_vector(15 downto 0);
    signal call14_1523 : std_logic_vector(15 downto 0);
    signal call15_1526 : std_logic_vector(15 downto 0);
    signal call16_1539 : std_logic_vector(15 downto 0);
    signal call18_1551 : std_logic_vector(15 downto 0);
    signal call1_1502 : std_logic_vector(15 downto 0);
    signal call20_1554 : std_logic_vector(15 downto 0);
    signal call22_1557 : std_logic_vector(15 downto 0);
    signal call3_1505 : std_logic_vector(15 downto 0);
    signal call5_1508 : std_logic_vector(15 downto 0);
    signal call7_1511 : std_logic_vector(15 downto 0);
    signal call9_1514 : std_logic_vector(15 downto 0);
    signal call_1499 : std_logic_vector(15 downto 0);
    signal cmp101_1781 : std_logic_vector(0 downto 0);
    signal cmp112_1806 : std_logic_vector(0 downto 0);
    signal cmp_1755 : std_logic_vector(0 downto 0);
    signal conv107_1801 : std_logic_vector(31 downto 0);
    signal conv110_1596 : std_logic_vector(31 downto 0);
    signal conv17_1543 : std_logic_vector(31 downto 0);
    signal conv61_1668 : std_logic_vector(63 downto 0);
    signal conv64_1584 : std_logic_vector(63 downto 0);
    signal conv66_1672 : std_logic_vector(63 downto 0);
    signal conv69_1588 : std_logic_vector(63 downto 0);
    signal conv71_1676 : std_logic_vector(63 downto 0);
    signal conv85_1744 : std_logic_vector(31 downto 0);
    signal conv89_1592 : std_logic_vector(31 downto 0);
    signal conv_1530 : std_logic_vector(31 downto 0);
    signal idxprom81_1729 : std_logic_vector(63 downto 0);
    signal idxprom_1706 : std_logic_vector(63 downto 0);
    signal inc105_1785 : std_logic_vector(15 downto 0);
    signal inc105x_xinput_dim0x_x2_1790 : std_logic_vector(15 downto 0);
    signal inc_1776 : std_logic_vector(15 downto 0);
    signal indvar_1605 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_1839 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_1827 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_1626 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_1821 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_1619 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_1797 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_1814 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1612 : std_logic_vector(15 downto 0);
    signal mul50_1659 : std_logic_vector(15 downto 0);
    signal mul72_1681 : std_logic_vector(63 downto 0);
    signal mul74_1691 : std_logic_vector(63 downto 0);
    signal mul_1649 : std_logic_vector(15 downto 0);
    signal ptr_deref_1716_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1716_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1716_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1716_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1716_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1738_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1738_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1738_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1738_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1738_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1738_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_1536 : std_logic_vector(31 downto 0);
    signal shr111126_1602 : std_logic_vector(31 downto 0);
    signal shr80_1723 : std_logic_vector(63 downto 0);
    signal shr_1702 : std_logic_vector(31 downto 0);
    signal sub44_1654 : std_logic_vector(15 downto 0);
    signal sub57_1580 : std_logic_vector(15 downto 0);
    signal sub58_1664 : std_logic_vector(15 downto 0);
    signal sub_1569 : std_logic_vector(15 downto 0);
    signal tmp1_1639 : std_logic_vector(31 downto 0);
    signal tmp78_1717 : std_logic_vector(63 downto 0);
    signal type_cast_1534_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1562_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1573_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1600_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1609_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1611_wire : std_logic_vector(31 downto 0);
    signal type_cast_1616_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1618_wire : std_logic_vector(15 downto 0);
    signal type_cast_1623_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1625_wire : std_logic_vector(15 downto 0);
    signal type_cast_1630_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1632_wire : std_logic_vector(15 downto 0);
    signal type_cast_1637_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1700_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1721_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1727_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1748_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1766_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1774_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1794_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1818_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1820_wire : std_logic_vector(15 downto 0);
    signal type_cast_1824_wire : std_logic_vector(15 downto 0);
    signal type_cast_1826_wire : std_logic_vector(15 downto 0);
    signal type_cast_1830_wire : std_logic_vector(15 downto 0);
    signal type_cast_1832_wire : std_logic_vector(15 downto 0);
    signal type_cast_1837_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1845_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_1711_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1711_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1711_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1711_resized_base_address <= "00000000000000";
    array_obj_ref_1734_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1734_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1734_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1734_resized_base_address <= "00000000000000";
    ptr_deref_1716_word_offset_0 <= "00000000000000";
    ptr_deref_1738_word_offset_0 <= "00000000000000";
    type_cast_1534_wire_constant <= "00000000000000000000000000010000";
    type_cast_1562_wire_constant <= "1111111111111111";
    type_cast_1573_wire_constant <= "1111111111111111";
    type_cast_1600_wire_constant <= "00000000000000000000000000000010";
    type_cast_1609_wire_constant <= "00000000000000000000000000000000";
    type_cast_1616_wire_constant <= "0000000000000000";
    type_cast_1623_wire_constant <= "0000000000000000";
    type_cast_1630_wire_constant <= "0000000000000000";
    type_cast_1637_wire_constant <= "00000000000000000000000000000100";
    type_cast_1700_wire_constant <= "00000000000000000000000000000010";
    type_cast_1721_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1727_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_1748_wire_constant <= "00000000000000000000000000000100";
    type_cast_1766_wire_constant <= "0000000000000100";
    type_cast_1774_wire_constant <= "0000000000000001";
    type_cast_1794_wire_constant <= "0000000000000000";
    type_cast_1818_wire_constant <= "0000000000000000";
    type_cast_1837_wire_constant <= "00000000000000000000000000000001";
    type_cast_1845_wire_constant <= "0000000000000001";
    phi_stmt_1605: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1609_wire_constant & type_cast_1611_wire;
      req <= phi_stmt_1605_req_0 & phi_stmt_1605_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1605",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1605_ack_0,
          idata => idata,
          odata => indvar_1605,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1605
    phi_stmt_1612: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1616_wire_constant & type_cast_1618_wire;
      req <= phi_stmt_1612_req_0 & phi_stmt_1612_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1612",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1612_ack_0,
          idata => idata,
          odata => input_dim2x_x1_1612,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1612
    phi_stmt_1619: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1623_wire_constant & type_cast_1625_wire;
      req <= phi_stmt_1619_req_0 & phi_stmt_1619_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1619",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1619_ack_0,
          idata => idata,
          odata => input_dim1x_x1_1619,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1619
    phi_stmt_1626: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1630_wire_constant & type_cast_1632_wire;
      req <= phi_stmt_1626_req_0 & phi_stmt_1626_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1626",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1626_ack_0,
          idata => idata,
          odata => input_dim0x_x2_1626,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1626
    phi_stmt_1814: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1818_wire_constant & type_cast_1820_wire;
      req <= phi_stmt_1814_req_0 & phi_stmt_1814_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1814",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1814_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_1814,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1814
    phi_stmt_1821: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1824_wire & type_cast_1826_wire;
      req <= phi_stmt_1821_req_0 & phi_stmt_1821_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1821",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1821_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_1821,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1821
    phi_stmt_1827: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1830_wire & type_cast_1832_wire;
      req <= phi_stmt_1827_req_0 & phi_stmt_1827_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1827",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1827_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_1827,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1827
    -- flow-through select operator MUX_1796_inst
    input_dim1x_x2_1797 <= type_cast_1794_wire_constant when (cmp101_1781(0) /=  '0') else inc_1776;
    addr_of_1712_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1712_final_reg_req_0;
      addr_of_1712_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1712_final_reg_req_1;
      addr_of_1712_final_reg_ack_1<= rack(0);
      addr_of_1712_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1712_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1711_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx77_1713,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1735_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1735_final_reg_req_0;
      addr_of_1735_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1735_final_reg_req_1;
      addr_of_1735_final_reg_ack_1<= rack(0);
      addr_of_1735_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1735_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1734_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx82_1736,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1529_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1529_inst_req_0;
      type_cast_1529_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1529_inst_req_1;
      type_cast_1529_inst_ack_1<= rack(0);
      type_cast_1529_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1529_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_1526,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1530,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1542_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1542_inst_req_0;
      type_cast_1542_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1542_inst_req_1;
      type_cast_1542_inst_ack_1<= rack(0);
      type_cast_1542_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1542_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_1539,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_1543,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1583_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1583_inst_req_0;
      type_cast_1583_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1583_inst_req_1;
      type_cast_1583_inst_ack_1<= rack(0);
      type_cast_1583_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1583_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_1557,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv64_1584,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1587_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1587_inst_req_0;
      type_cast_1587_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1587_inst_req_1;
      type_cast_1587_inst_ack_1<= rack(0);
      type_cast_1587_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1587_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_1554,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv69_1588,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1591_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1591_inst_req_0;
      type_cast_1591_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1591_inst_req_1;
      type_cast_1591_inst_ack_1<= rack(0);
      type_cast_1591_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1591_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_1505,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv89_1592,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1595_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1595_inst_req_0;
      type_cast_1595_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1595_inst_req_1;
      type_cast_1595_inst_ack_1<= rack(0);
      type_cast_1595_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1595_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1499,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv110_1596,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1611_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1611_inst_req_0;
      type_cast_1611_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1611_inst_req_1;
      type_cast_1611_inst_ack_1<= rack(0);
      type_cast_1611_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1611_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1839,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1611_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1618_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1618_inst_req_0;
      type_cast_1618_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1618_inst_req_1;
      type_cast_1618_inst_ack_1<= rack(0);
      type_cast_1618_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1618_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_1814,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1618_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1625_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1625_inst_req_0;
      type_cast_1625_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1625_inst_req_1;
      type_cast_1625_inst_ack_1<= rack(0);
      type_cast_1625_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1625_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_1821,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1625_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1632_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1632_inst_req_0;
      type_cast_1632_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1632_inst_req_1;
      type_cast_1632_inst_ack_1<= rack(0);
      type_cast_1632_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1632_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_1827,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1632_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1667_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1667_inst_req_0;
      type_cast_1667_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1667_inst_req_1;
      type_cast_1667_inst_ack_1<= rack(0);
      type_cast_1667_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1667_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1612,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv61_1668,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1671_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1671_inst_req_0;
      type_cast_1671_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1671_inst_req_1;
      type_cast_1671_inst_ack_1<= rack(0);
      type_cast_1671_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1671_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub58_1664,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv66_1672,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1675_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1675_inst_req_0;
      type_cast_1675_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1675_inst_req_1;
      type_cast_1675_inst_ack_1<= rack(0);
      type_cast_1675_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1675_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub44_1654,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv71_1676,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1705_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1705_inst_req_0;
      type_cast_1705_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1705_inst_req_1;
      type_cast_1705_inst_ack_1<= rack(0);
      type_cast_1705_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1705_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr_1702,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_1706,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1743_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1743_inst_req_0;
      type_cast_1743_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1743_inst_req_1;
      type_cast_1743_inst_ack_1<= rack(0);
      type_cast_1743_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1743_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1612,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv85_1744,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1784_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1784_inst_req_0;
      type_cast_1784_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1784_inst_req_1;
      type_cast_1784_inst_ack_1<= rack(0);
      type_cast_1784_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1784_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp101_1781,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc105_1785,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1800_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1800_inst_req_0;
      type_cast_1800_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1800_inst_req_1;
      type_cast_1800_inst_ack_1<= rack(0);
      type_cast_1800_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1800_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc105x_xinput_dim0x_x2_1790,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv107_1801,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1820_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1820_inst_req_0;
      type_cast_1820_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1820_inst_req_1;
      type_cast_1820_inst_ack_1<= rack(0);
      type_cast_1820_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1820_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add93_1768,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1820_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1824_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1824_inst_req_0;
      type_cast_1824_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1824_inst_req_1;
      type_cast_1824_inst_ack_1<= rack(0);
      type_cast_1824_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1824_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_1619,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1824_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1826_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1826_inst_req_0;
      type_cast_1826_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1826_inst_req_1;
      type_cast_1826_inst_ack_1<= rack(0);
      type_cast_1826_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1826_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_1797,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1826_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1830_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1830_inst_req_0;
      type_cast_1830_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1830_inst_req_1;
      type_cast_1830_inst_ack_1<= rack(0);
      type_cast_1830_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1830_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc105x_xinput_dim0x_x2_1790,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1830_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1832_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1832_inst_req_0;
      type_cast_1832_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1832_inst_req_1;
      type_cast_1832_inst_ack_1<= rack(0);
      type_cast_1832_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1832_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_1626,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1832_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1711_index_1_rename
    process(R_idxprom_1710_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_1710_resized;
      ov(13 downto 0) := iv;
      R_idxprom_1710_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1711_index_1_resize
    process(idxprom_1706) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_1706;
      ov := iv(13 downto 0);
      R_idxprom_1710_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1711_root_address_inst
    process(array_obj_ref_1711_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1711_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1711_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1734_index_1_rename
    process(R_idxprom81_1733_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom81_1733_resized;
      ov(13 downto 0) := iv;
      R_idxprom81_1733_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1734_index_1_resize
    process(idxprom81_1729) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom81_1729;
      ov := iv(13 downto 0);
      R_idxprom81_1733_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1734_root_address_inst
    process(array_obj_ref_1734_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1734_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1734_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1716_addr_0
    process(ptr_deref_1716_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1716_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1716_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1716_base_resize
    process(arrayidx77_1713) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx77_1713;
      ov := iv(13 downto 0);
      ptr_deref_1716_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1716_gather_scatter
    process(ptr_deref_1716_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1716_data_0;
      ov(63 downto 0) := iv;
      tmp78_1717 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1716_root_address_inst
    process(ptr_deref_1716_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1716_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1716_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1738_addr_0
    process(ptr_deref_1738_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1738_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1738_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1738_base_resize
    process(arrayidx82_1736) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx82_1736;
      ov := iv(13 downto 0);
      ptr_deref_1738_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1738_gather_scatter
    process(tmp78_1717) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp78_1717;
      ov(63 downto 0) := iv;
      ptr_deref_1738_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1738_root_address_inst
    process(ptr_deref_1738_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1738_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1738_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1756_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_1755;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1756_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1756_branch_req_0,
          ack0 => if_stmt_1756_branch_ack_0,
          ack1 => if_stmt_1756_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1807_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp112_1806;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1807_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1807_branch_req_0,
          ack0 => if_stmt_1807_branch_ack_0,
          ack1 => if_stmt_1807_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1563_inst
    process(call7_1511) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_1511, type_cast_1562_wire_constant, tmp_var);
      add41_1564 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1574_inst
    process(call9_1514) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_1514, type_cast_1573_wire_constant, tmp_var);
      add54_1575 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1653_inst
    process(sub_1569, mul_1649) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_1569, mul_1649, tmp_var);
      sub44_1654 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1663_inst
    process(sub57_1580, mul50_1659) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub57_1580, mul50_1659, tmp_var);
      sub58_1664 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1767_inst
    process(input_dim2x_x1_1612) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_1612, type_cast_1766_wire_constant, tmp_var);
      add93_1768 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1775_inst
    process(input_dim1x_x1_1619) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_1619, type_cast_1774_wire_constant, tmp_var);
      inc_1776 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1789_inst
    process(inc105_1785, input_dim0x_x2_1626) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc105_1785, input_dim0x_x2_1626, tmp_var);
      inc105x_xinput_dim0x_x2_1790 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1643_inst
    process(add_1548, tmp1_1639) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_1548, tmp1_1639, tmp_var);
      add_src_0x_x0_1644 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1749_inst
    process(conv85_1744) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv85_1744, type_cast_1748_wire_constant, tmp_var);
      add86_1750 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1838_inst
    process(indvar_1605) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1605, type_cast_1837_wire_constant, tmp_var);
      indvarx_xnext_1839 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1685_inst
    process(mul72_1681, conv66_1672) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul72_1681, conv66_1672, tmp_var);
      add73_1686 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1695_inst
    process(mul74_1691, conv61_1668) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul74_1691, conv61_1668, tmp_var);
      add75_1696 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1728_inst
    process(shr80_1723) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr80_1723, type_cast_1727_wire_constant, tmp_var);
      idxprom81_1729 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1780_inst
    process(inc_1776, call1_1502) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_1776, call1_1502, tmp_var);
      cmp101_1781 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1805_inst
    process(conv107_1801, shr111126_1602) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv107_1801, shr111126_1602, tmp_var);
      cmp112_1806 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1601_inst
    process(conv110_1596) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv110_1596, type_cast_1600_wire_constant, tmp_var);
      shr111126_1602 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1701_inst
    process(add_src_0x_x0_1644) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_1644, type_cast_1700_wire_constant, tmp_var);
      shr_1702 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1722_inst
    process(add75_1696) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add75_1696, type_cast_1721_wire_constant, tmp_var);
      shr80_1723 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1648_inst
    process(input_dim0x_x2_1626, call13_1520) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x2_1626, call13_1520, tmp_var);
      mul_1649 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1658_inst
    process(input_dim1x_x1_1619, call13_1520) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_1619, call13_1520, tmp_var);
      mul50_1659 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1638_inst
    process(indvar_1605) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_1605, type_cast_1637_wire_constant, tmp_var);
      tmp1_1639 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1680_inst
    process(conv71_1676, conv69_1588) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv71_1676, conv69_1588, tmp_var);
      mul72_1681 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1690_inst
    process(add73_1686, conv64_1584) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add73_1686, conv64_1584, tmp_var);
      mul74_1691 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1547_inst
    process(shl_1536, conv17_1543) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_1536, conv17_1543, tmp_var);
      add_1548 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1535_inst
    process(conv_1530) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_1530, type_cast_1534_wire_constant, tmp_var);
      shl_1536 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1568_inst
    process(add41_1564, call14_1523) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add41_1564, call14_1523, tmp_var);
      sub_1569 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1579_inst
    process(add54_1575, call14_1523) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add54_1575, call14_1523, tmp_var);
      sub57_1580 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1754_inst
    process(add86_1750, conv89_1592) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add86_1750, conv89_1592, tmp_var);
      cmp_1755 <= tmp_var; --
    end process;
    -- shared split operator group (28) : array_obj_ref_1711_index_offset 
    ApIntAdd_group_28: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_1710_scaled;
      array_obj_ref_1711_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1711_index_offset_req_0;
      array_obj_ref_1711_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1711_index_offset_req_1;
      array_obj_ref_1711_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_28_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_28_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : array_obj_ref_1734_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom81_1733_scaled;
      array_obj_ref_1734_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1734_index_offset_req_0;
      array_obj_ref_1734_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1734_index_offset_req_1;
      array_obj_ref_1734_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared load operator group (0) : ptr_deref_1716_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1716_load_0_req_0;
      ptr_deref_1716_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1716_load_0_req_1;
      ptr_deref_1716_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1716_word_address_0;
      ptr_deref_1716_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_1738_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1738_store_0_req_0;
      ptr_deref_1738_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1738_store_0_req_1;
      ptr_deref_1738_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1738_word_address_0;
      data_in <= ptr_deref_1738_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block0_start_1516_inst RPIPE_Block0_start_1525_inst RPIPE_Block0_start_1522_inst RPIPE_Block0_start_1538_inst RPIPE_Block0_start_1519_inst RPIPE_Block0_start_1513_inst RPIPE_Block0_start_1510_inst RPIPE_Block0_start_1553_inst RPIPE_Block0_start_1550_inst RPIPE_Block0_start_1498_inst RPIPE_Block0_start_1501_inst RPIPE_Block0_start_1556_inst RPIPE_Block0_start_1507_inst RPIPE_Block0_start_1504_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block0_start_1516_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block0_start_1525_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block0_start_1522_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block0_start_1538_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block0_start_1519_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block0_start_1513_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block0_start_1510_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block0_start_1553_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block0_start_1550_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block0_start_1498_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block0_start_1501_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block0_start_1556_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block0_start_1507_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block0_start_1504_inst_req_0;
      RPIPE_Block0_start_1516_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block0_start_1525_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block0_start_1522_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block0_start_1538_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block0_start_1519_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block0_start_1513_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block0_start_1510_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block0_start_1553_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block0_start_1550_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block0_start_1498_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block0_start_1501_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block0_start_1556_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block0_start_1507_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block0_start_1504_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block0_start_1516_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block0_start_1525_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block0_start_1522_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block0_start_1538_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block0_start_1519_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block0_start_1513_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block0_start_1510_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block0_start_1553_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block0_start_1550_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block0_start_1498_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block0_start_1501_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block0_start_1556_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block0_start_1507_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block0_start_1504_inst_req_1;
      RPIPE_Block0_start_1516_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block0_start_1525_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block0_start_1522_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block0_start_1538_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block0_start_1519_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block0_start_1513_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block0_start_1510_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block0_start_1553_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block0_start_1550_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block0_start_1498_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block0_start_1501_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block0_start_1556_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block0_start_1507_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block0_start_1504_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call11_1517 <= data_out(223 downto 208);
      call15_1526 <= data_out(207 downto 192);
      call14_1523 <= data_out(191 downto 176);
      call16_1539 <= data_out(175 downto 160);
      call13_1520 <= data_out(159 downto 144);
      call9_1514 <= data_out(143 downto 128);
      call7_1511 <= data_out(127 downto 112);
      call20_1554 <= data_out(111 downto 96);
      call18_1551 <= data_out(95 downto 80);
      call_1499 <= data_out(79 downto 64);
      call1_1502 <= data_out(63 downto 48);
      call22_1557 <= data_out(47 downto 32);
      call5_1508 <= data_out(31 downto 16);
      call3_1505 <= data_out(15 downto 0);
      Block0_start_read_0_gI: SplitGuardInterface generic map(name => "Block0_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_start_read_0: InputPortRevised -- 
        generic map ( name => "Block0_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_start_pipe_read_req(0),
          oack => Block0_start_pipe_read_ack(0),
          odata => Block0_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block0_done_1843_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block0_done_1843_inst_req_0;
      WPIPE_Block0_done_1843_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block0_done_1843_inst_req_1;
      WPIPE_Block0_done_1843_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_1845_wire_constant;
      Block0_done_write_0_gI: SplitGuardInterface generic map(name => "Block0_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_done_pipe_write_req(0),
          oack => Block0_done_pipe_write_ack(0),
          odata => Block0_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeA_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeB is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeB;
architecture convTransposeB_arch of convTransposeB is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeB_CP_4772_start: Boolean;
  signal convTransposeB_CP_4772_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_1885_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1878_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1875_inst_ack_0 : boolean;
  signal type_cast_1898_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1878_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1854_inst_ack_0 : boolean;
  signal type_cast_2185_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1875_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1906_inst_req_1 : boolean;
  signal type_cast_1898_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1875_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1875_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1857_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1866_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1857_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1866_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1860_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1857_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1860_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1854_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1854_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1854_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1866_inst_req_1 : boolean;
  signal type_cast_2187_inst_req_0 : boolean;
  signal type_cast_2187_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1909_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1909_inst_ack_1 : boolean;
  signal phi_stmt_1967_ack_0 : boolean;
  signal RPIPE_Block1_start_1906_inst_ack_0 : boolean;
  signal phi_stmt_2182_req_1 : boolean;
  signal type_cast_2185_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1881_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1872_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1881_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1872_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1906_inst_ack_1 : boolean;
  signal type_cast_1898_inst_req_0 : boolean;
  signal type_cast_1973_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1878_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1878_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1912_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1912_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1912_inst_ack_1 : boolean;
  signal type_cast_1945_inst_req_0 : boolean;
  signal type_cast_1945_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1909_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1909_inst_ack_0 : boolean;
  signal type_cast_1898_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1872_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1881_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1872_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1881_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1894_inst_ack_1 : boolean;
  signal phi_stmt_1967_req_1 : boolean;
  signal RPIPE_Block1_start_1894_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1860_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1906_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1866_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1860_inst_req_0 : boolean;
  signal type_cast_1957_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1894_inst_ack_0 : boolean;
  signal type_cast_1957_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1894_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1869_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1869_inst_req_1 : boolean;
  signal type_cast_1953_inst_req_1 : boolean;
  signal type_cast_1953_inst_ack_1 : boolean;
  signal type_cast_2187_inst_req_1 : boolean;
  signal type_cast_1953_inst_req_0 : boolean;
  signal type_cast_1953_inst_ack_0 : boolean;
  signal type_cast_2187_inst_ack_1 : boolean;
  signal type_cast_1973_inst_req_1 : boolean;
  signal type_cast_1885_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1869_inst_ack_0 : boolean;
  signal type_cast_1949_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1863_inst_ack_1 : boolean;
  signal type_cast_1885_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1869_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1863_inst_req_1 : boolean;
  signal type_cast_1957_inst_req_1 : boolean;
  signal type_cast_1957_inst_ack_1 : boolean;
  signal type_cast_1885_inst_ack_0 : boolean;
  signal type_cast_1949_inst_ack_1 : boolean;
  signal type_cast_1949_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1863_inst_ack_0 : boolean;
  signal type_cast_1949_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1863_inst_req_0 : boolean;
  signal type_cast_2028_inst_req_0 : boolean;
  signal type_cast_1945_inst_req_1 : boolean;
  signal type_cast_1945_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1857_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1912_inst_req_1 : boolean;
  signal phi_stmt_1974_ack_0 : boolean;
  signal type_cast_2028_inst_ack_0 : boolean;
  signal type_cast_2028_inst_req_1 : boolean;
  signal type_cast_2028_inst_ack_1 : boolean;
  signal type_cast_2032_inst_req_0 : boolean;
  signal type_cast_2032_inst_ack_0 : boolean;
  signal type_cast_2032_inst_req_1 : boolean;
  signal type_cast_2032_inst_ack_1 : boolean;
  signal type_cast_2036_inst_req_0 : boolean;
  signal type_cast_2036_inst_ack_0 : boolean;
  signal type_cast_2036_inst_req_1 : boolean;
  signal type_cast_2036_inst_ack_1 : boolean;
  signal type_cast_2066_inst_req_0 : boolean;
  signal type_cast_2066_inst_ack_0 : boolean;
  signal type_cast_2066_inst_req_1 : boolean;
  signal type_cast_2066_inst_ack_1 : boolean;
  signal phi_stmt_2188_req_0 : boolean;
  signal type_cast_2191_inst_ack_1 : boolean;
  signal type_cast_2191_inst_req_1 : boolean;
  signal array_obj_ref_2072_index_offset_req_0 : boolean;
  signal array_obj_ref_2072_index_offset_ack_0 : boolean;
  signal array_obj_ref_2072_index_offset_req_1 : boolean;
  signal array_obj_ref_2072_index_offset_ack_1 : boolean;
  signal addr_of_2073_final_reg_req_0 : boolean;
  signal addr_of_2073_final_reg_ack_0 : boolean;
  signal phi_stmt_2188_ack_0 : boolean;
  signal addr_of_2073_final_reg_req_1 : boolean;
  signal addr_of_2073_final_reg_ack_1 : boolean;
  signal type_cast_2191_inst_ack_0 : boolean;
  signal type_cast_2191_inst_req_0 : boolean;
  signal phi_stmt_2182_ack_0 : boolean;
  signal ptr_deref_2077_load_0_req_0 : boolean;
  signal ptr_deref_2077_load_0_ack_0 : boolean;
  signal phi_stmt_2175_ack_0 : boolean;
  signal ptr_deref_2077_load_0_req_1 : boolean;
  signal ptr_deref_2077_load_0_ack_1 : boolean;
  signal array_obj_ref_2095_index_offset_req_0 : boolean;
  signal array_obj_ref_2095_index_offset_ack_0 : boolean;
  signal array_obj_ref_2095_index_offset_req_1 : boolean;
  signal array_obj_ref_2095_index_offset_ack_1 : boolean;
  signal addr_of_2096_final_reg_req_0 : boolean;
  signal addr_of_2096_final_reg_ack_0 : boolean;
  signal phi_stmt_2175_req_0 : boolean;
  signal addr_of_2096_final_reg_req_1 : boolean;
  signal addr_of_2096_final_reg_ack_1 : boolean;
  signal type_cast_2178_inst_ack_1 : boolean;
  signal ptr_deref_2099_store_0_req_0 : boolean;
  signal ptr_deref_2099_store_0_ack_0 : boolean;
  signal type_cast_2178_inst_req_1 : boolean;
  signal phi_stmt_2188_req_1 : boolean;
  signal ptr_deref_2099_store_0_req_1 : boolean;
  signal phi_stmt_2175_req_1 : boolean;
  signal ptr_deref_2099_store_0_ack_1 : boolean;
  signal type_cast_2104_inst_req_0 : boolean;
  signal type_cast_2104_inst_ack_0 : boolean;
  signal type_cast_2104_inst_req_1 : boolean;
  signal type_cast_2104_inst_ack_1 : boolean;
  signal if_stmt_2117_branch_req_0 : boolean;
  signal if_stmt_2117_branch_ack_1 : boolean;
  signal type_cast_2178_inst_ack_0 : boolean;
  signal if_stmt_2117_branch_ack_0 : boolean;
  signal type_cast_2178_inst_req_0 : boolean;
  signal type_cast_2193_inst_ack_1 : boolean;
  signal type_cast_2145_inst_req_0 : boolean;
  signal type_cast_2145_inst_ack_0 : boolean;
  signal type_cast_2145_inst_req_1 : boolean;
  signal type_cast_2145_inst_ack_1 : boolean;
  signal type_cast_2161_inst_req_0 : boolean;
  signal type_cast_2161_inst_ack_0 : boolean;
  signal type_cast_2161_inst_req_1 : boolean;
  signal type_cast_2161_inst_ack_1 : boolean;
  signal if_stmt_2168_branch_req_0 : boolean;
  signal if_stmt_2168_branch_ack_1 : boolean;
  signal if_stmt_2168_branch_ack_0 : boolean;
  signal phi_stmt_1988_ack_0 : boolean;
  signal phi_stmt_1981_ack_0 : boolean;
  signal type_cast_2193_inst_req_1 : boolean;
  signal WPIPE_Block1_done_2204_inst_req_0 : boolean;
  signal WPIPE_Block1_done_2204_inst_ack_0 : boolean;
  signal WPIPE_Block1_done_2204_inst_req_1 : boolean;
  signal WPIPE_Block1_done_2204_inst_ack_1 : boolean;
  signal type_cast_1991_inst_req_0 : boolean;
  signal type_cast_1991_inst_ack_0 : boolean;
  signal type_cast_1991_inst_req_1 : boolean;
  signal phi_stmt_2182_req_0 : boolean;
  signal type_cast_1991_inst_ack_1 : boolean;
  signal phi_stmt_1988_req_0 : boolean;
  signal phi_stmt_1981_req_0 : boolean;
  signal type_cast_1973_inst_ack_0 : boolean;
  signal phi_stmt_1974_req_0 : boolean;
  signal phi_stmt_1967_req_0 : boolean;
  signal type_cast_2193_inst_ack_0 : boolean;
  signal type_cast_1993_inst_req_0 : boolean;
  signal type_cast_1993_inst_ack_0 : boolean;
  signal type_cast_2185_inst_ack_1 : boolean;
  signal type_cast_1993_inst_req_1 : boolean;
  signal type_cast_2185_inst_req_1 : boolean;
  signal type_cast_1993_inst_ack_1 : boolean;
  signal phi_stmt_1988_req_1 : boolean;
  signal type_cast_2193_inst_req_0 : boolean;
  signal type_cast_1987_inst_req_0 : boolean;
  signal type_cast_1987_inst_ack_0 : boolean;
  signal type_cast_1987_inst_req_1 : boolean;
  signal type_cast_1987_inst_ack_1 : boolean;
  signal phi_stmt_1981_req_1 : boolean;
  signal type_cast_1973_inst_req_0 : boolean;
  signal type_cast_1980_inst_req_0 : boolean;
  signal type_cast_1980_inst_ack_0 : boolean;
  signal type_cast_1980_inst_req_1 : boolean;
  signal type_cast_1980_inst_ack_1 : boolean;
  signal phi_stmt_1974_req_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeB_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeB_CP_4772_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeB_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_4772_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeB_CP_4772_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_4772_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeB_CP_4772: Block -- control-path 
    signal convTransposeB_CP_4772_elements: BooleanArray(127 downto 0);
    -- 
  begin -- 
    convTransposeB_CP_4772_elements(0) <= convTransposeB_CP_4772_start;
    convTransposeB_CP_4772_symbol <= convTransposeB_CP_4772_elements(78);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 branch_block_stmt_1852/branch_block_stmt_1852__entry__
      -- CP-element group 0: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913__entry__
      -- CP-element group 0: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/$entry
      -- CP-element group 0: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/type_cast_1898_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1854_sample_start_
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1854_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/type_cast_1885_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1854_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1852/$entry
      -- CP-element group 0: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/type_cast_1885_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/type_cast_1898_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/type_cast_1898_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/type_cast_1885_Update/cr
      -- 
    rr_4820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(0), ack => RPIPE_Block1_start_1854_inst_req_0); -- 
    cr_4993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(0), ack => type_cast_1898_inst_req_1); -- 
    cr_4965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(0), ack => type_cast_1885_inst_req_1); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	127 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	86 
    -- CP-element group 1: 	87 
    -- CP-element group 1: 	89 
    -- CP-element group 1: 	90 
    -- CP-element group 1: 	92 
    -- CP-element group 1: 	93 
    -- CP-element group 1: 	95 
    -- CP-element group 1: 	96 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_1852/merge_stmt_2174__exit__
      -- CP-element group 1: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_1852/assign_stmt_2200__exit__
      -- CP-element group 1: 	 branch_block_stmt_1852/assign_stmt_2200__entry__
      -- CP-element group 1: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/type_cast_1973/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1852/assign_stmt_2200/$entry
      -- CP-element group 1: 	 branch_block_stmt_1852/assign_stmt_2200/$exit
      -- CP-element group 1: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/type_cast_1973/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1988/$entry
      -- CP-element group 1: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1988/phi_stmt_1988_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1988/phi_stmt_1988_sources/type_cast_1993/$entry
      -- CP-element group 1: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1988/phi_stmt_1988_sources/type_cast_1993/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1988/phi_stmt_1988_sources/type_cast_1993/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1988/phi_stmt_1988_sources/type_cast_1993/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1988/phi_stmt_1988_sources/type_cast_1993/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1988/phi_stmt_1988_sources/type_cast_1993/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1981/$entry
      -- CP-element group 1: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1981/phi_stmt_1981_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1981/phi_stmt_1981_sources/type_cast_1987/$entry
      -- CP-element group 1: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1981/phi_stmt_1981_sources/type_cast_1987/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1981/phi_stmt_1981_sources/type_cast_1987/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1981/phi_stmt_1981_sources/type_cast_1987/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1981/phi_stmt_1981_sources/type_cast_1987/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1981/phi_stmt_1981_sources/type_cast_1987/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/type_cast_1973/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1974/$entry
      -- CP-element group 1: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1974/phi_stmt_1974_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1974/phi_stmt_1974_sources/type_cast_1980/$entry
      -- CP-element group 1: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1974/phi_stmt_1974_sources/type_cast_1980/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1974/phi_stmt_1974_sources/type_cast_1980/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1974/phi_stmt_1974_sources/type_cast_1980/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1974/phi_stmt_1974_sources/type_cast_1980/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1974/phi_stmt_1974_sources/type_cast_1980/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1967/$entry
      -- CP-element group 1: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/type_cast_1973/$entry
      -- CP-element group 1: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/type_cast_1973/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/type_cast_1973/SplitProtocol/Sample/$entry
      -- 
    cr_5595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(1), ack => type_cast_1973_inst_req_1); -- 
    rr_5521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(1), ack => type_cast_1993_inst_req_0); -- 
    cr_5526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(1), ack => type_cast_1993_inst_req_1); -- 
    rr_5544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(1), ack => type_cast_1987_inst_req_0); -- 
    cr_5549_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5549_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(1), ack => type_cast_1987_inst_req_1); -- 
    rr_5590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(1), ack => type_cast_1973_inst_req_0); -- 
    rr_5567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(1), ack => type_cast_1980_inst_req_0); -- 
    cr_5572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(1), ack => type_cast_1980_inst_req_1); -- 
    convTransposeB_CP_4772_elements(1) <= convTransposeB_CP_4772_elements(127);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1854_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1854_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1854_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1854_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1854_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1854_Update/cr
      -- 
    ra_4821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1854_inst_ack_0, ack => convTransposeB_CP_4772_elements(2)); -- 
    cr_4825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(2), ack => RPIPE_Block1_start_1854_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1857_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1854_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1854_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1854_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1857_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1857_sample_start_
      -- 
    ca_4826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1854_inst_ack_1, ack => convTransposeB_CP_4772_elements(3)); -- 
    rr_4834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(3), ack => RPIPE_Block1_start_1857_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1857_Update/cr
      -- CP-element group 4: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1857_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1857_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1857_update_start_
      -- CP-element group 4: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1857_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1857_Sample/ra
      -- 
    ra_4835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1857_inst_ack_0, ack => convTransposeB_CP_4772_elements(4)); -- 
    cr_4839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(4), ack => RPIPE_Block1_start_1857_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1857_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1857_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1860_Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1860_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1857_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1860_sample_start_
      -- 
    ca_4840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1857_inst_ack_1, ack => convTransposeB_CP_4772_elements(5)); -- 
    rr_4848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(5), ack => RPIPE_Block1_start_1860_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1860_Update/cr
      -- CP-element group 6: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1860_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1860_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1860_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1860_update_start_
      -- CP-element group 6: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1860_sample_completed_
      -- 
    ra_4849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1860_inst_ack_0, ack => convTransposeB_CP_4772_elements(6)); -- 
    cr_4853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(6), ack => RPIPE_Block1_start_1860_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1863_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1863_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1860_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1860_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1860_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1863_Sample/rr
      -- 
    ca_4854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1860_inst_ack_1, ack => convTransposeB_CP_4772_elements(7)); -- 
    rr_4862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(7), ack => RPIPE_Block1_start_1863_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1863_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1863_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1863_update_start_
      -- CP-element group 8: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1863_Update/cr
      -- CP-element group 8: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1863_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1863_Sample/ra
      -- 
    ra_4863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1863_inst_ack_0, ack => convTransposeB_CP_4772_elements(8)); -- 
    cr_4867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(8), ack => RPIPE_Block1_start_1863_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1866_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1866_Sample/rr
      -- CP-element group 9: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1863_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1866_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1863_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1863_Update/$exit
      -- 
    ca_4868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1863_inst_ack_1, ack => convTransposeB_CP_4772_elements(9)); -- 
    rr_4876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(9), ack => RPIPE_Block1_start_1866_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1866_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1866_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1866_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1866_update_start_
      -- CP-element group 10: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1866_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1866_Update/$entry
      -- 
    ra_4877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1866_inst_ack_0, ack => convTransposeB_CP_4772_elements(10)); -- 
    cr_4881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(10), ack => RPIPE_Block1_start_1866_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1866_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1866_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1869_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1866_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1869_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1869_Sample/$entry
      -- 
    ca_4882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1866_inst_ack_1, ack => convTransposeB_CP_4772_elements(11)); -- 
    rr_4890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(11), ack => RPIPE_Block1_start_1869_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1869_update_start_
      -- CP-element group 12: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1869_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1869_Update/cr
      -- CP-element group 12: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1869_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1869_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1869_Sample/$exit
      -- 
    ra_4891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1869_inst_ack_0, ack => convTransposeB_CP_4772_elements(12)); -- 
    cr_4895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(12), ack => RPIPE_Block1_start_1869_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1872_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1869_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1872_Sample/rr
      -- CP-element group 13: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1872_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1869_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1869_Update/$exit
      -- 
    ca_4896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1869_inst_ack_1, ack => convTransposeB_CP_4772_elements(13)); -- 
    rr_4904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(13), ack => RPIPE_Block1_start_1872_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1872_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1872_Update/cr
      -- CP-element group 14: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1872_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1872_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1872_update_start_
      -- CP-element group 14: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1872_sample_completed_
      -- 
    ra_4905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1872_inst_ack_0, ack => convTransposeB_CP_4772_elements(14)); -- 
    cr_4909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(14), ack => RPIPE_Block1_start_1872_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1875_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1875_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1875_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1872_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1872_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1872_update_completed_
      -- 
    ca_4910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1872_inst_ack_1, ack => convTransposeB_CP_4772_elements(15)); -- 
    rr_4918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(15), ack => RPIPE_Block1_start_1875_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1875_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1875_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1875_Update/cr
      -- CP-element group 16: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1875_update_start_
      -- CP-element group 16: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1875_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1875_Update/$entry
      -- 
    ra_4919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1875_inst_ack_0, ack => convTransposeB_CP_4772_elements(16)); -- 
    cr_4923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(16), ack => RPIPE_Block1_start_1875_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1878_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1875_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1875_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1878_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1878_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1875_Update/$exit
      -- 
    ca_4924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1875_inst_ack_1, ack => convTransposeB_CP_4772_elements(17)); -- 
    rr_4932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(17), ack => RPIPE_Block1_start_1878_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1878_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1878_Update/cr
      -- CP-element group 18: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1878_update_start_
      -- CP-element group 18: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1878_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1878_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1878_Update/$entry
      -- 
    ra_4933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1878_inst_ack_0, ack => convTransposeB_CP_4772_elements(18)); -- 
    cr_4937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(18), ack => RPIPE_Block1_start_1878_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1878_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1881_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1878_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1881_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1881_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1878_Update/$exit
      -- 
    ca_4938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1878_inst_ack_1, ack => convTransposeB_CP_4772_elements(19)); -- 
    rr_4946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(19), ack => RPIPE_Block1_start_1881_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1881_Update/cr
      -- CP-element group 20: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1881_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1881_update_start_
      -- CP-element group 20: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1881_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1881_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1881_Sample/$exit
      -- 
    ra_4947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1881_inst_ack_0, ack => convTransposeB_CP_4772_elements(20)); -- 
    cr_4951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(20), ack => RPIPE_Block1_start_1881_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/type_cast_1885_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/type_cast_1885_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1881_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/type_cast_1885_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1881_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1881_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1894_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1894_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1894_sample_start_
      -- 
    ca_4952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1881_inst_ack_1, ack => convTransposeB_CP_4772_elements(21)); -- 
    rr_4960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(21), ack => type_cast_1885_inst_req_0); -- 
    rr_4974_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4974_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(21), ack => RPIPE_Block1_start_1894_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/type_cast_1885_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/type_cast_1885_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/type_cast_1885_Sample/ra
      -- 
    ra_4961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1885_inst_ack_0, ack => convTransposeB_CP_4772_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/type_cast_1885_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/type_cast_1885_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/type_cast_1885_Update/$exit
      -- 
    ca_4966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1885_inst_ack_1, ack => convTransposeB_CP_4772_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1894_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1894_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1894_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1894_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1894_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1894_sample_completed_
      -- 
    ra_4975_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1894_inst_ack_0, ack => convTransposeB_CP_4772_elements(24)); -- 
    cr_4979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(24), ack => RPIPE_Block1_start_1894_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/type_cast_1898_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1906_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/type_cast_1898_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/type_cast_1898_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1906_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1894_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1894_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1906_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1894_update_completed_
      -- 
    ca_4980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1894_inst_ack_1, ack => convTransposeB_CP_4772_elements(25)); -- 
    rr_4988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(25), ack => type_cast_1898_inst_req_0); -- 
    rr_5002_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5002_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(25), ack => RPIPE_Block1_start_1906_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/type_cast_1898_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/type_cast_1898_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/type_cast_1898_sample_completed_
      -- 
    ra_4989_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1898_inst_ack_0, ack => convTransposeB_CP_4772_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/type_cast_1898_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/type_cast_1898_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/type_cast_1898_update_completed_
      -- 
    ca_4994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1898_inst_ack_1, ack => convTransposeB_CP_4772_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1906_Update/cr
      -- CP-element group 28: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1906_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1906_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1906_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1906_update_start_
      -- CP-element group 28: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1906_Update/$entry
      -- 
    ra_5003_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1906_inst_ack_0, ack => convTransposeB_CP_4772_elements(28)); -- 
    cr_5007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(28), ack => RPIPE_Block1_start_1906_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1909_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1906_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1906_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1909_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1909_Sample/rr
      -- CP-element group 29: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1906_Update/$exit
      -- 
    ca_5008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1906_inst_ack_1, ack => convTransposeB_CP_4772_elements(29)); -- 
    rr_5016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(29), ack => RPIPE_Block1_start_1909_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1909_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1909_Update/cr
      -- CP-element group 30: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1909_update_start_
      -- CP-element group 30: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1909_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1909_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1909_sample_completed_
      -- 
    ra_5017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1909_inst_ack_0, ack => convTransposeB_CP_4772_elements(30)); -- 
    cr_5021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(30), ack => RPIPE_Block1_start_1909_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1912_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1909_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1912_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1909_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1909_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1912_Sample/rr
      -- 
    ca_5022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1909_inst_ack_1, ack => convTransposeB_CP_4772_elements(31)); -- 
    rr_5030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(31), ack => RPIPE_Block1_start_1912_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1912_update_start_
      -- CP-element group 32: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1912_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1912_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1912_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1912_Update/cr
      -- CP-element group 32: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1912_Update/$entry
      -- 
    ra_5031_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1912_inst_ack_0, ack => convTransposeB_CP_4772_elements(32)); -- 
    cr_5035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(32), ack => RPIPE_Block1_start_1912_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1912_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1912_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/RPIPE_Block1_start_1912_Update/$exit
      -- 
    ca_5036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1912_inst_ack_1, ack => convTransposeB_CP_4772_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34: 	41 
    -- CP-element group 34: 	42 
    -- CP-element group 34:  members (28) 
      -- CP-element group 34: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913/$exit
      -- CP-element group 34: 	 branch_block_stmt_1852/assign_stmt_1855_to_assign_stmt_1913__exit__
      -- CP-element group 34: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964__entry__
      -- CP-element group 34: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1949_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1945_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1945_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1945_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/$entry
      -- CP-element group 34: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1945_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1945_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1957_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1957_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1957_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1957_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1957_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1953_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1953_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1953_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1953_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1949_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1949_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1953_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1953_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1957_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1949_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1949_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1945_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1949_update_start_
      -- 
    rr_5047_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5047_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(34), ack => type_cast_1945_inst_req_0); -- 
    rr_5089_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5089_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(34), ack => type_cast_1957_inst_req_0); -- 
    cr_5080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(34), ack => type_cast_1953_inst_req_1); -- 
    rr_5075_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5075_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(34), ack => type_cast_1953_inst_req_0); -- 
    rr_5061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(34), ack => type_cast_1949_inst_req_0); -- 
    cr_5094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(34), ack => type_cast_1957_inst_req_1); -- 
    cr_5066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(34), ack => type_cast_1949_inst_req_1); -- 
    cr_5052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(34), ack => type_cast_1945_inst_req_1); -- 
    convTransposeB_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(23) & convTransposeB_CP_4772_elements(27) & convTransposeB_CP_4772_elements(33);
      gj_convTransposeB_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1945_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1945_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1945_sample_completed_
      -- 
    ra_5048_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1945_inst_ack_0, ack => convTransposeB_CP_4772_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	43 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1945_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1945_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1945_Update/ca
      -- 
    ca_5053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1945_inst_ack_1, ack => convTransposeB_CP_4772_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1949_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1949_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1949_Sample/ra
      -- 
    ra_5062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1949_inst_ack_0, ack => convTransposeB_CP_4772_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	43 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1949_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1949_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1949_update_completed_
      -- 
    ca_5067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1949_inst_ack_1, ack => convTransposeB_CP_4772_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1953_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1953_Sample/ra
      -- CP-element group 39: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1953_sample_completed_
      -- 
    ra_5076_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1953_inst_ack_0, ack => convTransposeB_CP_4772_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	43 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1953_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1953_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1953_update_completed_
      -- 
    ca_5081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1953_inst_ack_1, ack => convTransposeB_CP_4772_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	34 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1957_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1957_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1957_sample_completed_
      -- 
    ra_5090_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1957_inst_ack_0, ack => convTransposeB_CP_4772_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	34 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1957_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1957_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/type_cast_1957_Update/ca
      -- 
    ca_5095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1957_inst_ack_1, ack => convTransposeB_CP_4772_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  place  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	36 
    -- CP-element group 43: 	38 
    -- CP-element group 43: 	40 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	79 
    -- CP-element group 43: 	80 
    -- CP-element group 43: 	82 
    -- CP-element group 43: 	83 
    -- CP-element group 43: 	84 
    -- CP-element group 43:  members (18) 
      -- CP-element group 43: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964__exit__
      -- CP-element group 43: 	 branch_block_stmt_1852/entry_whilex_xbody
      -- CP-element group 43: 	 branch_block_stmt_1852/assign_stmt_1920_to_assign_stmt_1964/$exit
      -- CP-element group 43: 	 branch_block_stmt_1852/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 43: 	 branch_block_stmt_1852/entry_whilex_xbody_PhiReq/phi_stmt_1988/$entry
      -- CP-element group 43: 	 branch_block_stmt_1852/entry_whilex_xbody_PhiReq/phi_stmt_1988/phi_stmt_1988_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1852/entry_whilex_xbody_PhiReq/phi_stmt_1988/phi_stmt_1988_sources/type_cast_1991/$entry
      -- CP-element group 43: 	 branch_block_stmt_1852/entry_whilex_xbody_PhiReq/phi_stmt_1988/phi_stmt_1988_sources/type_cast_1991/SplitProtocol/$entry
      -- CP-element group 43: 	 branch_block_stmt_1852/entry_whilex_xbody_PhiReq/phi_stmt_1988/phi_stmt_1988_sources/type_cast_1991/SplitProtocol/Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_1852/entry_whilex_xbody_PhiReq/phi_stmt_1988/phi_stmt_1988_sources/type_cast_1991/SplitProtocol/Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_1852/entry_whilex_xbody_PhiReq/phi_stmt_1988/phi_stmt_1988_sources/type_cast_1991/SplitProtocol/Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_1852/entry_whilex_xbody_PhiReq/phi_stmt_1988/phi_stmt_1988_sources/type_cast_1991/SplitProtocol/Update/cr
      -- CP-element group 43: 	 branch_block_stmt_1852/entry_whilex_xbody_PhiReq/phi_stmt_1981/$entry
      -- CP-element group 43: 	 branch_block_stmt_1852/entry_whilex_xbody_PhiReq/phi_stmt_1981/phi_stmt_1981_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1852/entry_whilex_xbody_PhiReq/phi_stmt_1974/$entry
      -- CP-element group 43: 	 branch_block_stmt_1852/entry_whilex_xbody_PhiReq/phi_stmt_1974/phi_stmt_1974_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1852/entry_whilex_xbody_PhiReq/phi_stmt_1967/$entry
      -- CP-element group 43: 	 branch_block_stmt_1852/entry_whilex_xbody_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/$entry
      -- 
    rr_5471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(43), ack => type_cast_1991_inst_req_0); -- 
    cr_5476_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5476_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(43), ack => type_cast_1991_inst_req_1); -- 
    convTransposeB_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(36) & convTransposeB_CP_4772_elements(38) & convTransposeB_CP_4772_elements(40) & convTransposeB_CP_4772_elements(42);
      gj_convTransposeB_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	104 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2028_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2028_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2028_Sample/ra
      -- 
    ra_5107_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2028_inst_ack_0, ack => convTransposeB_CP_4772_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	104 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	58 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2028_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2028_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2028_Update/ca
      -- 
    ca_5112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2028_inst_ack_1, ack => convTransposeB_CP_4772_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	104 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2032_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2032_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2032_Sample/ra
      -- 
    ra_5121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2032_inst_ack_0, ack => convTransposeB_CP_4772_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	104 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	58 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2032_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2032_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2032_Update/ca
      -- 
    ca_5126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2032_inst_ack_1, ack => convTransposeB_CP_4772_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	104 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2036_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2036_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2036_Sample/ra
      -- 
    ra_5135_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2036_inst_ack_0, ack => convTransposeB_CP_4772_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	104 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2036_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2036_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2036_Update/ca
      -- 
    ca_5140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2036_inst_ack_1, ack => convTransposeB_CP_4772_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	104 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2066_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2066_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2066_Sample/ra
      -- 
    ra_5149_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2066_inst_ack_0, ack => convTransposeB_CP_4772_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	104 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (16) 
      -- CP-element group 51: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2066_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2066_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2066_Update/ca
      -- CP-element group 51: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2072_index_resized_1
      -- CP-element group 51: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2072_index_scaled_1
      -- CP-element group 51: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2072_index_computed_1
      -- CP-element group 51: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2072_index_resize_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2072_index_resize_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2072_index_resize_1/index_resize_req
      -- CP-element group 51: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2072_index_resize_1/index_resize_ack
      -- CP-element group 51: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2072_index_scale_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2072_index_scale_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2072_index_scale_1/scale_rename_req
      -- CP-element group 51: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2072_index_scale_1/scale_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2072_final_index_sum_regn_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2072_final_index_sum_regn_Sample/req
      -- 
    ca_5154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2066_inst_ack_1, ack => convTransposeB_CP_4772_elements(51)); -- 
    req_5179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(51), ack => array_obj_ref_2072_index_offset_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	68 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2072_final_index_sum_regn_sample_complete
      -- CP-element group 52: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2072_final_index_sum_regn_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2072_final_index_sum_regn_Sample/ack
      -- 
    ack_5180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2072_index_offset_ack_0, ack => convTransposeB_CP_4772_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	104 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (11) 
      -- CP-element group 53: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/addr_of_2073_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2072_root_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2072_offset_calculated
      -- CP-element group 53: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2072_final_index_sum_regn_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2072_final_index_sum_regn_Update/ack
      -- CP-element group 53: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2072_base_plus_offset/$entry
      -- CP-element group 53: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2072_base_plus_offset/$exit
      -- CP-element group 53: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2072_base_plus_offset/sum_rename_req
      -- CP-element group 53: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2072_base_plus_offset/sum_rename_ack
      -- CP-element group 53: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/addr_of_2073_request/$entry
      -- CP-element group 53: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/addr_of_2073_request/req
      -- 
    ack_5185_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2072_index_offset_ack_1, ack => convTransposeB_CP_4772_elements(53)); -- 
    req_5194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(53), ack => addr_of_2073_final_reg_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/addr_of_2073_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/addr_of_2073_request/$exit
      -- CP-element group 54: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/addr_of_2073_request/ack
      -- 
    ack_5195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2073_final_reg_ack_0, ack => convTransposeB_CP_4772_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	104 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (24) 
      -- CP-element group 55: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/addr_of_2073_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/addr_of_2073_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/addr_of_2073_complete/ack
      -- CP-element group 55: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2077_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2077_base_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2077_word_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2077_root_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2077_base_address_resized
      -- CP-element group 55: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2077_base_addr_resize/$entry
      -- CP-element group 55: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2077_base_addr_resize/$exit
      -- CP-element group 55: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2077_base_addr_resize/base_resize_req
      -- CP-element group 55: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2077_base_addr_resize/base_resize_ack
      -- CP-element group 55: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2077_base_plus_offset/$entry
      -- CP-element group 55: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2077_base_plus_offset/$exit
      -- CP-element group 55: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2077_base_plus_offset/sum_rename_req
      -- CP-element group 55: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2077_base_plus_offset/sum_rename_ack
      -- CP-element group 55: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2077_word_addrgen/$entry
      -- CP-element group 55: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2077_word_addrgen/$exit
      -- CP-element group 55: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2077_word_addrgen/root_register_req
      -- CP-element group 55: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2077_word_addrgen/root_register_ack
      -- CP-element group 55: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2077_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2077_Sample/word_access_start/$entry
      -- CP-element group 55: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2077_Sample/word_access_start/word_0/$entry
      -- CP-element group 55: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2077_Sample/word_access_start/word_0/rr
      -- 
    ack_5200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2073_final_reg_ack_1, ack => convTransposeB_CP_4772_elements(55)); -- 
    rr_5233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(55), ack => ptr_deref_2077_load_0_req_0); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (5) 
      -- CP-element group 56: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2077_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2077_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2077_Sample/word_access_start/$exit
      -- CP-element group 56: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2077_Sample/word_access_start/word_0/$exit
      -- CP-element group 56: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2077_Sample/word_access_start/word_0/ra
      -- 
    ra_5234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2077_load_0_ack_0, ack => convTransposeB_CP_4772_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	104 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (9) 
      -- CP-element group 57: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2077_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2077_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2077_Update/word_access_complete/$exit
      -- CP-element group 57: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2077_Update/word_access_complete/word_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2077_Update/word_access_complete/word_0/ca
      -- CP-element group 57: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2077_Update/ptr_deref_2077_Merge/$entry
      -- CP-element group 57: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2077_Update/ptr_deref_2077_Merge/$exit
      -- CP-element group 57: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2077_Update/ptr_deref_2077_Merge/merge_req
      -- CP-element group 57: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2077_Update/ptr_deref_2077_Merge/merge_ack
      -- 
    ca_5245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2077_load_0_ack_1, ack => convTransposeB_CP_4772_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	45 
    -- CP-element group 58: 	47 
    -- CP-element group 58: 	49 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (13) 
      -- CP-element group 58: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2095_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2095_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2095_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2095_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2095_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2095_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2095_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2095_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2095_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2095_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2095_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2095_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2095_final_index_sum_regn_Sample/req
      -- 
    req_5275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(58), ack => array_obj_ref_2095_index_offset_req_0); -- 
    convTransposeB_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(45) & convTransposeB_CP_4772_elements(47) & convTransposeB_CP_4772_elements(49);
      gj_convTransposeB_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	68 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2095_final_index_sum_regn_sample_complete
      -- CP-element group 59: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2095_final_index_sum_regn_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2095_final_index_sum_regn_Sample/ack
      -- 
    ack_5276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2095_index_offset_ack_0, ack => convTransposeB_CP_4772_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	104 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (11) 
      -- CP-element group 60: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/addr_of_2096_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2095_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2095_offset_calculated
      -- CP-element group 60: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2095_final_index_sum_regn_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2095_final_index_sum_regn_Update/ack
      -- CP-element group 60: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2095_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2095_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2095_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2095_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/addr_of_2096_request/$entry
      -- CP-element group 60: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/addr_of_2096_request/req
      -- 
    ack_5281_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2095_index_offset_ack_1, ack => convTransposeB_CP_4772_elements(60)); -- 
    req_5290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(60), ack => addr_of_2096_final_reg_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/addr_of_2096_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/addr_of_2096_request/$exit
      -- CP-element group 61: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/addr_of_2096_request/ack
      -- 
    ack_5291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2096_final_reg_ack_0, ack => convTransposeB_CP_4772_elements(61)); -- 
    -- CP-element group 62:  fork  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	104 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (19) 
      -- CP-element group 62: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/addr_of_2096_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/addr_of_2096_complete/$exit
      -- CP-element group 62: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/addr_of_2096_complete/ack
      -- CP-element group 62: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2099_base_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2099_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2099_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2099_base_address_resized
      -- CP-element group 62: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2099_base_addr_resize/$entry
      -- CP-element group 62: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2099_base_addr_resize/$exit
      -- CP-element group 62: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2099_base_addr_resize/base_resize_req
      -- CP-element group 62: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2099_base_addr_resize/base_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2099_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2099_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2099_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2099_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2099_word_addrgen/$entry
      -- CP-element group 62: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2099_word_addrgen/$exit
      -- CP-element group 62: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2099_word_addrgen/root_register_req
      -- CP-element group 62: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2099_word_addrgen/root_register_ack
      -- 
    ack_5296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2096_final_reg_ack_1, ack => convTransposeB_CP_4772_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2099_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2099_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2099_Sample/ptr_deref_2099_Split/$entry
      -- CP-element group 63: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2099_Sample/ptr_deref_2099_Split/$exit
      -- CP-element group 63: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2099_Sample/ptr_deref_2099_Split/split_req
      -- CP-element group 63: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2099_Sample/ptr_deref_2099_Split/split_ack
      -- CP-element group 63: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2099_Sample/word_access_start/$entry
      -- CP-element group 63: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2099_Sample/word_access_start/word_0/$entry
      -- CP-element group 63: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2099_Sample/word_access_start/word_0/rr
      -- 
    rr_5334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(63), ack => ptr_deref_2099_store_0_req_0); -- 
    convTransposeB_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(57) & convTransposeB_CP_4772_elements(62);
      gj_convTransposeB_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2099_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2099_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2099_Sample/word_access_start/$exit
      -- CP-element group 64: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2099_Sample/word_access_start/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2099_Sample/word_access_start/word_0/ra
      -- 
    ra_5335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2099_store_0_ack_0, ack => convTransposeB_CP_4772_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	104 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	68 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2099_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2099_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2099_Update/word_access_complete/$exit
      -- CP-element group 65: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2099_Update/word_access_complete/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2099_Update/word_access_complete/word_0/ca
      -- 
    ca_5346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2099_store_0_ack_1, ack => convTransposeB_CP_4772_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	104 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2104_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2104_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2104_Sample/ra
      -- 
    ra_5355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2104_inst_ack_0, ack => convTransposeB_CP_4772_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	104 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2104_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2104_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2104_Update/ca
      -- 
    ca_5360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2104_inst_ack_1, ack => convTransposeB_CP_4772_elements(67)); -- 
    -- CP-element group 68:  branch  join  transition  place  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	52 
    -- CP-element group 68: 	59 
    -- CP-element group 68: 	65 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (10) 
      -- CP-element group 68: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116__exit__
      -- CP-element group 68: 	 branch_block_stmt_1852/if_stmt_2117__entry__
      -- CP-element group 68: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/$exit
      -- CP-element group 68: 	 branch_block_stmt_1852/if_stmt_2117_dead_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1852/if_stmt_2117_eval_test/$entry
      -- CP-element group 68: 	 branch_block_stmt_1852/if_stmt_2117_eval_test/$exit
      -- CP-element group 68: 	 branch_block_stmt_1852/if_stmt_2117_eval_test/branch_req
      -- CP-element group 68: 	 branch_block_stmt_1852/R_cmp_2118_place
      -- CP-element group 68: 	 branch_block_stmt_1852/if_stmt_2117_if_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1852/if_stmt_2117_else_link/$entry
      -- 
    branch_req_5368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(68), ack => if_stmt_2117_branch_req_0); -- 
    convTransposeB_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(52) & convTransposeB_CP_4772_elements(59) & convTransposeB_CP_4772_elements(65) & convTransposeB_CP_4772_elements(67);
      gj_convTransposeB_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	113 
    -- CP-element group 69: 	114 
    -- CP-element group 69: 	116 
    -- CP-element group 69: 	117 
    -- CP-element group 69: 	119 
    -- CP-element group 69: 	120 
    -- CP-element group 69:  members (40) 
      -- CP-element group 69: 	 branch_block_stmt_1852/assign_stmt_2129__entry__
      -- CP-element group 69: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2175/$entry
      -- CP-element group 69: 	 branch_block_stmt_1852/assign_stmt_2129__exit__
      -- CP-element group 69: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128
      -- CP-element group 69: 	 branch_block_stmt_1852/merge_stmt_2123__exit__
      -- CP-element group 69: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2187/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2187/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2187/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2187/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2187/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2187/$entry
      -- CP-element group 69: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2182/$entry
      -- CP-element group 69: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2191/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2191/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2191/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2191/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2191/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2191/$entry
      -- CP-element group 69: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2188/$entry
      -- CP-element group 69: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/type_cast_2178/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1852/merge_stmt_2123_PhiReqMerge
      -- CP-element group 69: 	 branch_block_stmt_1852/merge_stmt_2123_PhiAck/dummy
      -- CP-element group 69: 	 branch_block_stmt_1852/merge_stmt_2123_PhiAck/$exit
      -- CP-element group 69: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/type_cast_2178/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1852/if_stmt_2117_if_link/$exit
      -- CP-element group 69: 	 branch_block_stmt_1852/merge_stmt_2123_PhiAck/$entry
      -- CP-element group 69: 	 branch_block_stmt_1852/if_stmt_2117_if_link/if_choice_transition
      -- CP-element group 69: 	 branch_block_stmt_1852/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 69: 	 branch_block_stmt_1852/whilex_xbody_ifx_xthen
      -- CP-element group 69: 	 branch_block_stmt_1852/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/type_cast_2178/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1852/assign_stmt_2129/$entry
      -- CP-element group 69: 	 branch_block_stmt_1852/assign_stmt_2129/$exit
      -- CP-element group 69: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/type_cast_2178/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/type_cast_2178/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/type_cast_2178/$entry
      -- 
    if_choice_transition_5373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2117_branch_ack_1, ack => convTransposeB_CP_4772_elements(69)); -- 
    rr_5728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(69), ack => type_cast_2187_inst_req_0); -- 
    cr_5733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(69), ack => type_cast_2187_inst_req_1); -- 
    cr_5710_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5710_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(69), ack => type_cast_2191_inst_req_1); -- 
    rr_5705_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5705_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(69), ack => type_cast_2191_inst_req_0); -- 
    cr_5756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(69), ack => type_cast_2178_inst_req_1); -- 
    rr_5751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(69), ack => type_cast_2178_inst_req_0); -- 
    -- CP-element group 70:  fork  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70: 	74 
    -- CP-element group 70:  members (21) 
      -- CP-element group 70: 	 branch_block_stmt_1852/merge_stmt_2131__exit__
      -- CP-element group 70: 	 branch_block_stmt_1852/assign_stmt_2137_to_assign_stmt_2167__entry__
      -- CP-element group 70: 	 branch_block_stmt_1852/merge_stmt_2131_PhiAck/dummy
      -- CP-element group 70: 	 branch_block_stmt_1852/merge_stmt_2131_PhiAck/$exit
      -- CP-element group 70: 	 branch_block_stmt_1852/merge_stmt_2131_PhiAck/$entry
      -- CP-element group 70: 	 branch_block_stmt_1852/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 70: 	 branch_block_stmt_1852/merge_stmt_2131_PhiReqMerge
      -- CP-element group 70: 	 branch_block_stmt_1852/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_1852/if_stmt_2117_else_link/$exit
      -- CP-element group 70: 	 branch_block_stmt_1852/if_stmt_2117_else_link/else_choice_transition
      -- CP-element group 70: 	 branch_block_stmt_1852/whilex_xbody_ifx_xelse
      -- CP-element group 70: 	 branch_block_stmt_1852/assign_stmt_2137_to_assign_stmt_2167/$entry
      -- CP-element group 70: 	 branch_block_stmt_1852/assign_stmt_2137_to_assign_stmt_2167/type_cast_2145_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_1852/assign_stmt_2137_to_assign_stmt_2167/type_cast_2145_update_start_
      -- CP-element group 70: 	 branch_block_stmt_1852/assign_stmt_2137_to_assign_stmt_2167/type_cast_2145_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_1852/assign_stmt_2137_to_assign_stmt_2167/type_cast_2145_Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_1852/assign_stmt_2137_to_assign_stmt_2167/type_cast_2145_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1852/assign_stmt_2137_to_assign_stmt_2167/type_cast_2145_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_1852/assign_stmt_2137_to_assign_stmt_2167/type_cast_2161_update_start_
      -- CP-element group 70: 	 branch_block_stmt_1852/assign_stmt_2137_to_assign_stmt_2167/type_cast_2161_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1852/assign_stmt_2137_to_assign_stmt_2167/type_cast_2161_Update/cr
      -- 
    else_choice_transition_5377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2117_branch_ack_0, ack => convTransposeB_CP_4772_elements(70)); -- 
    rr_5393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(70), ack => type_cast_2145_inst_req_0); -- 
    cr_5398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(70), ack => type_cast_2145_inst_req_1); -- 
    cr_5412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(70), ack => type_cast_2161_inst_req_1); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_1852/assign_stmt_2137_to_assign_stmt_2167/type_cast_2145_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_1852/assign_stmt_2137_to_assign_stmt_2167/type_cast_2145_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_1852/assign_stmt_2137_to_assign_stmt_2167/type_cast_2145_Sample/ra
      -- 
    ra_5394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2145_inst_ack_0, ack => convTransposeB_CP_4772_elements(71)); -- 
    -- CP-element group 72:  transition  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (6) 
      -- CP-element group 72: 	 branch_block_stmt_1852/assign_stmt_2137_to_assign_stmt_2167/type_cast_2145_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_1852/assign_stmt_2137_to_assign_stmt_2167/type_cast_2145_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_1852/assign_stmt_2137_to_assign_stmt_2167/type_cast_2145_Update/ca
      -- CP-element group 72: 	 branch_block_stmt_1852/assign_stmt_2137_to_assign_stmt_2167/type_cast_2161_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_1852/assign_stmt_2137_to_assign_stmt_2167/type_cast_2161_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_1852/assign_stmt_2137_to_assign_stmt_2167/type_cast_2161_Sample/rr
      -- 
    ca_5399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2145_inst_ack_1, ack => convTransposeB_CP_4772_elements(72)); -- 
    rr_5407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(72), ack => type_cast_2161_inst_req_0); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1852/assign_stmt_2137_to_assign_stmt_2167/type_cast_2161_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_1852/assign_stmt_2137_to_assign_stmt_2167/type_cast_2161_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_1852/assign_stmt_2137_to_assign_stmt_2167/type_cast_2161_Sample/ra
      -- 
    ra_5408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2161_inst_ack_0, ack => convTransposeB_CP_4772_elements(73)); -- 
    -- CP-element group 74:  branch  transition  place  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	70 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (13) 
      -- CP-element group 74: 	 branch_block_stmt_1852/assign_stmt_2137_to_assign_stmt_2167__exit__
      -- CP-element group 74: 	 branch_block_stmt_1852/if_stmt_2168__entry__
      -- CP-element group 74: 	 branch_block_stmt_1852/assign_stmt_2137_to_assign_stmt_2167/$exit
      -- CP-element group 74: 	 branch_block_stmt_1852/assign_stmt_2137_to_assign_stmt_2167/type_cast_2161_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_1852/assign_stmt_2137_to_assign_stmt_2167/type_cast_2161_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_1852/assign_stmt_2137_to_assign_stmt_2167/type_cast_2161_Update/ca
      -- CP-element group 74: 	 branch_block_stmt_1852/if_stmt_2168_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1852/if_stmt_2168_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_1852/if_stmt_2168_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_1852/if_stmt_2168_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_1852/R_cmp117_2169_place
      -- CP-element group 74: 	 branch_block_stmt_1852/if_stmt_2168_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1852/if_stmt_2168_else_link/$entry
      -- 
    ca_5413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2161_inst_ack_1, ack => convTransposeB_CP_4772_elements(74)); -- 
    branch_req_5421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(74), ack => if_stmt_2168_branch_req_0); -- 
    -- CP-element group 75:  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (15) 
      -- CP-element group 75: 	 branch_block_stmt_1852/assign_stmt_2207__entry__
      -- CP-element group 75: 	 branch_block_stmt_1852/merge_stmt_2202__exit__
      -- CP-element group 75: 	 branch_block_stmt_1852/merge_stmt_2202_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_1852/merge_stmt_2202_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_1852/merge_stmt_2202_PhiAck/dummy
      -- CP-element group 75: 	 branch_block_stmt_1852/merge_stmt_2202_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_1852/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_1852/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_1852/if_stmt_2168_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_1852/if_stmt_2168_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_1852/ifx_xelse_whilex_xend
      -- CP-element group 75: 	 branch_block_stmt_1852/assign_stmt_2207/$entry
      -- CP-element group 75: 	 branch_block_stmt_1852/assign_stmt_2207/WPIPE_Block1_done_2204_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_1852/assign_stmt_2207/WPIPE_Block1_done_2204_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_1852/assign_stmt_2207/WPIPE_Block1_done_2204_Sample/req
      -- 
    if_choice_transition_5426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2168_branch_ack_1, ack => convTransposeB_CP_4772_elements(75)); -- 
    req_5446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(75), ack => WPIPE_Block1_done_2204_inst_req_0); -- 
    -- CP-element group 76:  fork  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	105 
    -- CP-element group 76: 	106 
    -- CP-element group 76: 	108 
    -- CP-element group 76: 	109 
    -- CP-element group 76: 	111 
    -- CP-element group 76:  members (22) 
      -- CP-element group 76: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2185/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2185/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2193/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2193/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2185/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2193/$entry
      -- CP-element group 76: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2185/$entry
      -- CP-element group 76: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2182/$entry
      -- CP-element group 76: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1852/if_stmt_2168_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_1852/if_stmt_2168_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128
      -- CP-element group 76: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2193/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2188/$entry
      -- CP-element group 76: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2193/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2175/$entry
      -- CP-element group 76: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2185/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2193/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2185/SplitProtocol/Update/$entry
      -- 
    else_choice_transition_5430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2168_branch_ack_0, ack => convTransposeB_CP_4772_elements(76)); -- 
    rr_5671_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5671_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(76), ack => type_cast_2185_inst_req_0); -- 
    cr_5653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(76), ack => type_cast_2193_inst_req_1); -- 
    cr_5676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(76), ack => type_cast_2185_inst_req_1); -- 
    rr_5648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(76), ack => type_cast_2193_inst_req_0); -- 
    -- CP-element group 77:  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (6) 
      -- CP-element group 77: 	 branch_block_stmt_1852/assign_stmt_2207/WPIPE_Block1_done_2204_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_1852/assign_stmt_2207/WPIPE_Block1_done_2204_update_start_
      -- CP-element group 77: 	 branch_block_stmt_1852/assign_stmt_2207/WPIPE_Block1_done_2204_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_1852/assign_stmt_2207/WPIPE_Block1_done_2204_Sample/ack
      -- CP-element group 77: 	 branch_block_stmt_1852/assign_stmt_2207/WPIPE_Block1_done_2204_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1852/assign_stmt_2207/WPIPE_Block1_done_2204_Update/req
      -- 
    ack_5447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2204_inst_ack_0, ack => convTransposeB_CP_4772_elements(77)); -- 
    req_5451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(77), ack => WPIPE_Block1_done_2204_inst_req_1); -- 
    -- CP-element group 78:  transition  place  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (16) 
      -- CP-element group 78: 	 branch_block_stmt_1852/merge_stmt_2209__exit__
      -- CP-element group 78: 	 branch_block_stmt_1852/branch_block_stmt_1852__exit__
      -- CP-element group 78: 	 branch_block_stmt_1852/return__
      -- CP-element group 78: 	 branch_block_stmt_1852/$exit
      -- CP-element group 78: 	 $exit
      -- CP-element group 78: 	 branch_block_stmt_1852/assign_stmt_2207__exit__
      -- CP-element group 78: 	 branch_block_stmt_1852/return___PhiReq/$entry
      -- CP-element group 78: 	 branch_block_stmt_1852/merge_stmt_2209_PhiReqMerge
      -- CP-element group 78: 	 branch_block_stmt_1852/assign_stmt_2207/$exit
      -- CP-element group 78: 	 branch_block_stmt_1852/assign_stmt_2207/WPIPE_Block1_done_2204_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_1852/assign_stmt_2207/WPIPE_Block1_done_2204_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_1852/assign_stmt_2207/WPIPE_Block1_done_2204_Update/ack
      -- CP-element group 78: 	 branch_block_stmt_1852/merge_stmt_2209_PhiAck/dummy
      -- CP-element group 78: 	 branch_block_stmt_1852/merge_stmt_2209_PhiAck/$exit
      -- CP-element group 78: 	 branch_block_stmt_1852/merge_stmt_2209_PhiAck/$entry
      -- CP-element group 78: 	 branch_block_stmt_1852/return___PhiReq/$exit
      -- 
    ack_5452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2204_inst_ack_1, ack => convTransposeB_CP_4772_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	43 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_1852/entry_whilex_xbody_PhiReq/phi_stmt_1988/phi_stmt_1988_sources/type_cast_1991/SplitProtocol/Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_1852/entry_whilex_xbody_PhiReq/phi_stmt_1988/phi_stmt_1988_sources/type_cast_1991/SplitProtocol/Sample/ra
      -- 
    ra_5472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1991_inst_ack_0, ack => convTransposeB_CP_4772_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	43 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_1852/entry_whilex_xbody_PhiReq/phi_stmt_1988/phi_stmt_1988_sources/type_cast_1991/SplitProtocol/Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_1852/entry_whilex_xbody_PhiReq/phi_stmt_1988/phi_stmt_1988_sources/type_cast_1991/SplitProtocol/Update/ca
      -- 
    ca_5477_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1991_inst_ack_1, ack => convTransposeB_CP_4772_elements(80)); -- 
    -- CP-element group 81:  join  transition  output  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	85 
    -- CP-element group 81:  members (5) 
      -- CP-element group 81: 	 branch_block_stmt_1852/entry_whilex_xbody_PhiReq/phi_stmt_1988/$exit
      -- CP-element group 81: 	 branch_block_stmt_1852/entry_whilex_xbody_PhiReq/phi_stmt_1988/phi_stmt_1988_sources/$exit
      -- CP-element group 81: 	 branch_block_stmt_1852/entry_whilex_xbody_PhiReq/phi_stmt_1988/phi_stmt_1988_sources/type_cast_1991/$exit
      -- CP-element group 81: 	 branch_block_stmt_1852/entry_whilex_xbody_PhiReq/phi_stmt_1988/phi_stmt_1988_sources/type_cast_1991/SplitProtocol/$exit
      -- CP-element group 81: 	 branch_block_stmt_1852/entry_whilex_xbody_PhiReq/phi_stmt_1988/phi_stmt_1988_req
      -- 
    phi_stmt_1988_req_5478_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1988_req_5478_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(81), ack => phi_stmt_1988_req_0); -- 
    convTransposeB_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(79) & convTransposeB_CP_4772_elements(80);
      gj_convTransposeB_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  transition  output  delay-element  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	43 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	85 
    -- CP-element group 82:  members (4) 
      -- CP-element group 82: 	 branch_block_stmt_1852/entry_whilex_xbody_PhiReq/phi_stmt_1981/$exit
      -- CP-element group 82: 	 branch_block_stmt_1852/entry_whilex_xbody_PhiReq/phi_stmt_1981/phi_stmt_1981_sources/$exit
      -- CP-element group 82: 	 branch_block_stmt_1852/entry_whilex_xbody_PhiReq/phi_stmt_1981/phi_stmt_1981_sources/type_cast_1985_konst_delay_trans
      -- CP-element group 82: 	 branch_block_stmt_1852/entry_whilex_xbody_PhiReq/phi_stmt_1981/phi_stmt_1981_req
      -- 
    phi_stmt_1981_req_5486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1981_req_5486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(82), ack => phi_stmt_1981_req_0); -- 
    -- Element group convTransposeB_CP_4772_elements(82) is a control-delay.
    cp_element_82_delay: control_delay_element  generic map(name => " 82_delay", delay_value => 1)  port map(req => convTransposeB_CP_4772_elements(43), ack => convTransposeB_CP_4772_elements(82), clk => clk, reset =>reset);
    -- CP-element group 83:  transition  output  delay-element  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	43 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (4) 
      -- CP-element group 83: 	 branch_block_stmt_1852/entry_whilex_xbody_PhiReq/phi_stmt_1974/$exit
      -- CP-element group 83: 	 branch_block_stmt_1852/entry_whilex_xbody_PhiReq/phi_stmt_1974/phi_stmt_1974_sources/$exit
      -- CP-element group 83: 	 branch_block_stmt_1852/entry_whilex_xbody_PhiReq/phi_stmt_1974/phi_stmt_1974_sources/type_cast_1978_konst_delay_trans
      -- CP-element group 83: 	 branch_block_stmt_1852/entry_whilex_xbody_PhiReq/phi_stmt_1974/phi_stmt_1974_req
      -- 
    phi_stmt_1974_req_5494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1974_req_5494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(83), ack => phi_stmt_1974_req_0); -- 
    -- Element group convTransposeB_CP_4772_elements(83) is a control-delay.
    cp_element_83_delay: control_delay_element  generic map(name => " 83_delay", delay_value => 1)  port map(req => convTransposeB_CP_4772_elements(43), ack => convTransposeB_CP_4772_elements(83), clk => clk, reset =>reset);
    -- CP-element group 84:  transition  output  delay-element  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	43 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (4) 
      -- CP-element group 84: 	 branch_block_stmt_1852/entry_whilex_xbody_PhiReq/phi_stmt_1967/$exit
      -- CP-element group 84: 	 branch_block_stmt_1852/entry_whilex_xbody_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/$exit
      -- CP-element group 84: 	 branch_block_stmt_1852/entry_whilex_xbody_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/type_cast_1971_konst_delay_trans
      -- CP-element group 84: 	 branch_block_stmt_1852/entry_whilex_xbody_PhiReq/phi_stmt_1967/phi_stmt_1967_req
      -- 
    phi_stmt_1967_req_5502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1967_req_5502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(84), ack => phi_stmt_1967_req_0); -- 
    -- Element group convTransposeB_CP_4772_elements(84) is a control-delay.
    cp_element_84_delay: control_delay_element  generic map(name => " 84_delay", delay_value => 1)  port map(req => convTransposeB_CP_4772_elements(43), ack => convTransposeB_CP_4772_elements(84), clk => clk, reset =>reset);
    -- CP-element group 85:  join  transition  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	81 
    -- CP-element group 85: 	82 
    -- CP-element group 85: 	83 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	99 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_1852/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(81) & convTransposeB_CP_4772_elements(82) & convTransposeB_CP_4772_elements(83) & convTransposeB_CP_4772_elements(84);
      gj_convTransposeB_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	1 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1988/phi_stmt_1988_sources/type_cast_1993/SplitProtocol/Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1988/phi_stmt_1988_sources/type_cast_1993/SplitProtocol/Sample/ra
      -- 
    ra_5522_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1993_inst_ack_0, ack => convTransposeB_CP_4772_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	1 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1988/phi_stmt_1988_sources/type_cast_1993/SplitProtocol/Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1988/phi_stmt_1988_sources/type_cast_1993/SplitProtocol/Update/ca
      -- 
    ca_5527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1993_inst_ack_1, ack => convTransposeB_CP_4772_elements(87)); -- 
    -- CP-element group 88:  join  transition  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	98 
    -- CP-element group 88:  members (5) 
      -- CP-element group 88: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1988/$exit
      -- CP-element group 88: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1988/phi_stmt_1988_sources/$exit
      -- CP-element group 88: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1988/phi_stmt_1988_sources/type_cast_1993/$exit
      -- CP-element group 88: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1988/phi_stmt_1988_sources/type_cast_1993/SplitProtocol/$exit
      -- CP-element group 88: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1988/phi_stmt_1988_req
      -- 
    phi_stmt_1988_req_5528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1988_req_5528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(88), ack => phi_stmt_1988_req_1); -- 
    convTransposeB_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(86) & convTransposeB_CP_4772_elements(87);
      gj_convTransposeB_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	1 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1981/phi_stmt_1981_sources/type_cast_1987/SplitProtocol/Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1981/phi_stmt_1981_sources/type_cast_1987/SplitProtocol/Sample/ra
      -- 
    ra_5545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1987_inst_ack_0, ack => convTransposeB_CP_4772_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	1 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1981/phi_stmt_1981_sources/type_cast_1987/SplitProtocol/Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1981/phi_stmt_1981_sources/type_cast_1987/SplitProtocol/Update/ca
      -- 
    ca_5550_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1987_inst_ack_1, ack => convTransposeB_CP_4772_elements(90)); -- 
    -- CP-element group 91:  join  transition  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	98 
    -- CP-element group 91:  members (5) 
      -- CP-element group 91: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1981/$exit
      -- CP-element group 91: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1981/phi_stmt_1981_sources/$exit
      -- CP-element group 91: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1981/phi_stmt_1981_sources/type_cast_1987/$exit
      -- CP-element group 91: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1981/phi_stmt_1981_sources/type_cast_1987/SplitProtocol/$exit
      -- CP-element group 91: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1981/phi_stmt_1981_req
      -- 
    phi_stmt_1981_req_5551_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1981_req_5551_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(91), ack => phi_stmt_1981_req_1); -- 
    convTransposeB_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(89) & convTransposeB_CP_4772_elements(90);
      gj_convTransposeB_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	1 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1974/phi_stmt_1974_sources/type_cast_1980/SplitProtocol/Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1974/phi_stmt_1974_sources/type_cast_1980/SplitProtocol/Sample/ra
      -- 
    ra_5568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1980_inst_ack_0, ack => convTransposeB_CP_4772_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	1 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1974/phi_stmt_1974_sources/type_cast_1980/SplitProtocol/Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1974/phi_stmt_1974_sources/type_cast_1980/SplitProtocol/Update/ca
      -- 
    ca_5573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1980_inst_ack_1, ack => convTransposeB_CP_4772_elements(93)); -- 
    -- CP-element group 94:  join  transition  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	98 
    -- CP-element group 94:  members (5) 
      -- CP-element group 94: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1974/$exit
      -- CP-element group 94: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1974/phi_stmt_1974_sources/$exit
      -- CP-element group 94: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1974/phi_stmt_1974_sources/type_cast_1980/$exit
      -- CP-element group 94: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1974/phi_stmt_1974_sources/type_cast_1980/SplitProtocol/$exit
      -- CP-element group 94: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1974/phi_stmt_1974_req
      -- 
    phi_stmt_1974_req_5574_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1974_req_5574_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(94), ack => phi_stmt_1974_req_1); -- 
    convTransposeB_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(92) & convTransposeB_CP_4772_elements(93);
      gj_convTransposeB_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	1 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/type_cast_1973/SplitProtocol/Sample/ra
      -- CP-element group 95: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/type_cast_1973/SplitProtocol/Sample/$exit
      -- 
    ra_5591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1973_inst_ack_0, ack => convTransposeB_CP_4772_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	1 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/type_cast_1973/SplitProtocol/Update/ca
      -- CP-element group 96: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/type_cast_1973/SplitProtocol/Update/$exit
      -- 
    ca_5596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1973_inst_ack_1, ack => convTransposeB_CP_4772_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1967/phi_stmt_1967_req
      -- CP-element group 97: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1967/$exit
      -- CP-element group 97: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/$exit
      -- CP-element group 97: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/type_cast_1973/$exit
      -- CP-element group 97: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/type_cast_1973/SplitProtocol/$exit
      -- 
    phi_stmt_1967_req_5597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1967_req_5597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(97), ack => phi_stmt_1967_req_1); -- 
    convTransposeB_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(95) & convTransposeB_CP_4772_elements(96);
      gj_convTransposeB_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	88 
    -- CP-element group 98: 	91 
    -- CP-element group 98: 	94 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_1852/ifx_xend128_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(88) & convTransposeB_CP_4772_elements(91) & convTransposeB_CP_4772_elements(94) & convTransposeB_CP_4772_elements(97);
      gj_convTransposeB_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  merge  fork  transition  place  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	85 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: 	101 
    -- CP-element group 99: 	102 
    -- CP-element group 99: 	103 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_1852/merge_stmt_1966_PhiAck/$entry
      -- CP-element group 99: 	 branch_block_stmt_1852/merge_stmt_1966_PhiReqMerge
      -- 
    convTransposeB_CP_4772_elements(99) <= OrReduce(convTransposeB_CP_4772_elements(85) & convTransposeB_CP_4772_elements(98));
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	104 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_1852/merge_stmt_1966_PhiAck/phi_stmt_1967_ack
      -- 
    phi_stmt_1967_ack_5602_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1967_ack_0, ack => convTransposeB_CP_4772_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	104 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_1852/merge_stmt_1966_PhiAck/phi_stmt_1974_ack
      -- 
    phi_stmt_1974_ack_5603_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1974_ack_0, ack => convTransposeB_CP_4772_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	99 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_1852/merge_stmt_1966_PhiAck/phi_stmt_1981_ack
      -- 
    phi_stmt_1981_ack_5604_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1981_ack_0, ack => convTransposeB_CP_4772_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	99 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_1852/merge_stmt_1966_PhiAck/phi_stmt_1988_ack
      -- 
    phi_stmt_1988_ack_5605_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1988_ack_0, ack => convTransposeB_CP_4772_elements(103)); -- 
    -- CP-element group 104:  join  fork  transition  place  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	100 
    -- CP-element group 104: 	101 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	44 
    -- CP-element group 104: 	45 
    -- CP-element group 104: 	46 
    -- CP-element group 104: 	47 
    -- CP-element group 104: 	48 
    -- CP-element group 104: 	49 
    -- CP-element group 104: 	50 
    -- CP-element group 104: 	51 
    -- CP-element group 104: 	53 
    -- CP-element group 104: 	55 
    -- CP-element group 104: 	57 
    -- CP-element group 104: 	60 
    -- CP-element group 104: 	62 
    -- CP-element group 104: 	65 
    -- CP-element group 104: 	66 
    -- CP-element group 104: 	67 
    -- CP-element group 104:  members (56) 
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116__entry__
      -- CP-element group 104: 	 branch_block_stmt_1852/merge_stmt_1966__exit__
      -- CP-element group 104: 	 branch_block_stmt_1852/merge_stmt_1966_PhiAck/$exit
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2028_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/$entry
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2028_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2028_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2028_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2028_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2028_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2032_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2032_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2032_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2032_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2032_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2032_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2036_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2036_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2036_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2036_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2036_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2036_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2066_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2066_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2066_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2066_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2066_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2066_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/addr_of_2073_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2072_final_index_sum_regn_update_start
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2072_final_index_sum_regn_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2072_final_index_sum_regn_Update/req
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/addr_of_2073_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/addr_of_2073_complete/req
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2077_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2077_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2077_Update/word_access_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2077_Update/word_access_complete/word_0/$entry
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2077_Update/word_access_complete/word_0/cr
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/addr_of_2096_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2095_final_index_sum_regn_update_start
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2095_final_index_sum_regn_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/array_obj_ref_2095_final_index_sum_regn_Update/req
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/addr_of_2096_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/addr_of_2096_complete/req
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2099_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2099_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2099_Update/word_access_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2099_Update/word_access_complete/word_0/$entry
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/ptr_deref_2099_Update/word_access_complete/word_0/cr
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2104_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2104_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2104_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2104_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2104_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1852/assign_stmt_2000_to_assign_stmt_2116/type_cast_2104_Update/cr
      -- 
    rr_5106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(104), ack => type_cast_2028_inst_req_0); -- 
    cr_5111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(104), ack => type_cast_2028_inst_req_1); -- 
    rr_5120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(104), ack => type_cast_2032_inst_req_0); -- 
    cr_5125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(104), ack => type_cast_2032_inst_req_1); -- 
    rr_5134_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5134_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(104), ack => type_cast_2036_inst_req_0); -- 
    cr_5139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(104), ack => type_cast_2036_inst_req_1); -- 
    rr_5148_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5148_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(104), ack => type_cast_2066_inst_req_0); -- 
    cr_5153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(104), ack => type_cast_2066_inst_req_1); -- 
    req_5184_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5184_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(104), ack => array_obj_ref_2072_index_offset_req_1); -- 
    req_5199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(104), ack => addr_of_2073_final_reg_req_1); -- 
    cr_5244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(104), ack => ptr_deref_2077_load_0_req_1); -- 
    req_5280_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5280_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(104), ack => array_obj_ref_2095_index_offset_req_1); -- 
    req_5295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(104), ack => addr_of_2096_final_reg_req_1); -- 
    cr_5345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(104), ack => ptr_deref_2099_store_0_req_1); -- 
    rr_5354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(104), ack => type_cast_2104_inst_req_0); -- 
    cr_5359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(104), ack => type_cast_2104_inst_req_1); -- 
    convTransposeB_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(100) & convTransposeB_CP_4772_elements(101) & convTransposeB_CP_4772_elements(102) & convTransposeB_CP_4772_elements(103);
      gj_convTransposeB_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	76 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2193/SplitProtocol/Sample/ra
      -- CP-element group 105: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2193/SplitProtocol/Sample/$exit
      -- 
    ra_5649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2193_inst_ack_0, ack => convTransposeB_CP_4772_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	76 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2193/SplitProtocol/Update/ca
      -- CP-element group 106: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2193/SplitProtocol/Update/$exit
      -- 
    ca_5654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2193_inst_ack_1, ack => convTransposeB_CP_4772_elements(106)); -- 
    -- CP-element group 107:  join  transition  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	112 
    -- CP-element group 107:  members (5) 
      -- CP-element group 107: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2193/SplitProtocol/$exit
      -- CP-element group 107: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2193/$exit
      -- CP-element group 107: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/$exit
      -- CP-element group 107: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2188/$exit
      -- CP-element group 107: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_req
      -- 
    phi_stmt_2188_req_5655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2188_req_5655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(107), ack => phi_stmt_2188_req_1); -- 
    convTransposeB_cp_element_group_107: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_107"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(105) & convTransposeB_CP_4772_elements(106);
      gj_convTransposeB_cp_element_group_107 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	76 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	110 
    -- CP-element group 108:  members (2) 
      -- CP-element group 108: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2185/SplitProtocol/Sample/ra
      -- CP-element group 108: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2185/SplitProtocol/Sample/$exit
      -- 
    ra_5672_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2185_inst_ack_0, ack => convTransposeB_CP_4772_elements(108)); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	76 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2185/SplitProtocol/Update/ca
      -- CP-element group 109: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2185/SplitProtocol/Update/$exit
      -- 
    ca_5677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2185_inst_ack_1, ack => convTransposeB_CP_4772_elements(109)); -- 
    -- CP-element group 110:  join  transition  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	108 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	112 
    -- CP-element group 110:  members (5) 
      -- CP-element group 110: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2185/SplitProtocol/$exit
      -- CP-element group 110: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2185/$exit
      -- CP-element group 110: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/$exit
      -- CP-element group 110: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2182/$exit
      -- CP-element group 110: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2182/phi_stmt_2182_req
      -- 
    phi_stmt_2182_req_5678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2182_req_5678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(110), ack => phi_stmt_2182_req_0); -- 
    convTransposeB_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(108) & convTransposeB_CP_4772_elements(109);
      gj_convTransposeB_cp_element_group_110 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  transition  output  delay-element  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	76 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (4) 
      -- CP-element group 111: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2175/phi_stmt_2175_req
      -- CP-element group 111: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/type_cast_2181_konst_delay_trans
      -- CP-element group 111: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/$exit
      -- CP-element group 111: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2175/$exit
      -- 
    phi_stmt_2175_req_5686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2175_req_5686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(111), ack => phi_stmt_2175_req_1); -- 
    -- Element group convTransposeB_CP_4772_elements(111) is a control-delay.
    cp_element_111_delay: control_delay_element  generic map(name => " 111_delay", delay_value => 1)  port map(req => convTransposeB_CP_4772_elements(76), ack => convTransposeB_CP_4772_elements(111), clk => clk, reset =>reset);
    -- CP-element group 112:  join  transition  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	107 
    -- CP-element group 112: 	110 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	123 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_1852/ifx_xelse_ifx_xend128_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(107) & convTransposeB_CP_4772_elements(110) & convTransposeB_CP_4772_elements(111);
      gj_convTransposeB_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	69 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2191/SplitProtocol/Sample/ra
      -- CP-element group 113: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2191/SplitProtocol/Sample/$exit
      -- 
    ra_5706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2191_inst_ack_0, ack => convTransposeB_CP_4772_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	69 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (2) 
      -- CP-element group 114: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2191/SplitProtocol/Update/ca
      -- CP-element group 114: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2191/SplitProtocol/Update/$exit
      -- 
    ca_5711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2191_inst_ack_1, ack => convTransposeB_CP_4772_elements(114)); -- 
    -- CP-element group 115:  join  transition  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	122 
    -- CP-element group 115:  members (5) 
      -- CP-element group 115: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_req
      -- CP-element group 115: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2191/SplitProtocol/$exit
      -- CP-element group 115: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2191/$exit
      -- CP-element group 115: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/$exit
      -- CP-element group 115: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2188/$exit
      -- 
    phi_stmt_2188_req_5712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2188_req_5712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(115), ack => phi_stmt_2188_req_0); -- 
    convTransposeB_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(113) & convTransposeB_CP_4772_elements(114);
      gj_convTransposeB_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	69 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (2) 
      -- CP-element group 116: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2187/SplitProtocol/Sample/ra
      -- CP-element group 116: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2187/SplitProtocol/Sample/$exit
      -- 
    ra_5729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2187_inst_ack_0, ack => convTransposeB_CP_4772_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	69 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2187/SplitProtocol/Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2187/SplitProtocol/Update/ca
      -- 
    ca_5734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2187_inst_ack_1, ack => convTransposeB_CP_4772_elements(117)); -- 
    -- CP-element group 118:  join  transition  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	122 
    -- CP-element group 118:  members (5) 
      -- CP-element group 118: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2182/phi_stmt_2182_req
      -- CP-element group 118: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2187/SplitProtocol/$exit
      -- CP-element group 118: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2187/$exit
      -- CP-element group 118: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/$exit
      -- CP-element group 118: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2182/$exit
      -- 
    phi_stmt_2182_req_5735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2182_req_5735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(118), ack => phi_stmt_2182_req_1); -- 
    convTransposeB_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(116) & convTransposeB_CP_4772_elements(117);
      gj_convTransposeB_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	69 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/type_cast_2178/SplitProtocol/Sample/ra
      -- CP-element group 119: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/type_cast_2178/SplitProtocol/Sample/$exit
      -- 
    ra_5752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2178_inst_ack_0, ack => convTransposeB_CP_4772_elements(119)); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	69 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/type_cast_2178/SplitProtocol/Update/ca
      -- CP-element group 120: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/type_cast_2178/SplitProtocol/Update/$exit
      -- 
    ca_5757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2178_inst_ack_1, ack => convTransposeB_CP_4772_elements(120)); -- 
    -- CP-element group 121:  join  transition  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (5) 
      -- CP-element group 121: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2175/$exit
      -- CP-element group 121: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2175/phi_stmt_2175_req
      -- CP-element group 121: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/type_cast_2178/SplitProtocol/$exit
      -- CP-element group 121: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/type_cast_2178/$exit
      -- CP-element group 121: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/$exit
      -- 
    phi_stmt_2175_req_5758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2175_req_5758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(121), ack => phi_stmt_2175_req_0); -- 
    convTransposeB_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(119) & convTransposeB_CP_4772_elements(120);
      gj_convTransposeB_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  join  transition  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	115 
    -- CP-element group 122: 	118 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_1852/ifx_xthen_ifx_xend128_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(115) & convTransposeB_CP_4772_elements(118) & convTransposeB_CP_4772_elements(121);
      gj_convTransposeB_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  merge  fork  transition  place  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	112 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123: 	125 
    -- CP-element group 123: 	126 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_1852/merge_stmt_2174_PhiReqMerge
      -- CP-element group 123: 	 branch_block_stmt_1852/merge_stmt_2174_PhiAck/$entry
      -- 
    convTransposeB_CP_4772_elements(123) <= OrReduce(convTransposeB_CP_4772_elements(112) & convTransposeB_CP_4772_elements(122));
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	127 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_1852/merge_stmt_2174_PhiAck/phi_stmt_2175_ack
      -- 
    phi_stmt_2175_ack_5763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2175_ack_0, ack => convTransposeB_CP_4772_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_1852/merge_stmt_2174_PhiAck/phi_stmt_2182_ack
      -- 
    phi_stmt_2182_ack_5764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2182_ack_0, ack => convTransposeB_CP_4772_elements(125)); -- 
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	123 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (1) 
      -- CP-element group 126: 	 branch_block_stmt_1852/merge_stmt_2174_PhiAck/phi_stmt_2188_ack
      -- 
    phi_stmt_2188_ack_5765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2188_ack_0, ack => convTransposeB_CP_4772_elements(126)); -- 
    -- CP-element group 127:  join  transition  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	124 
    -- CP-element group 127: 	125 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	1 
    -- CP-element group 127:  members (1) 
      -- CP-element group 127: 	 branch_block_stmt_1852/merge_stmt_2174_PhiAck/$exit
      -- 
    convTransposeB_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(124) & convTransposeB_CP_4772_elements(125) & convTransposeB_CP_4772_elements(126);
      gj_convTransposeB_cp_element_group_127 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(127), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom86_2094_resized : std_logic_vector(13 downto 0);
    signal R_idxprom86_2094_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2071_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2071_scaled : std_logic_vector(13 downto 0);
    signal add45_1926 : std_logic_vector(15 downto 0);
    signal add58_1937 : std_logic_vector(15 downto 0);
    signal add77_2047 : std_logic_vector(63 downto 0);
    signal add79_2057 : std_logic_vector(63 downto 0);
    signal add91_2111 : std_logic_vector(31 downto 0);
    signal add98_2129 : std_logic_vector(15 downto 0);
    signal add_1904 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_2005 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2072_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2072_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2072_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2072_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2072_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2072_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2095_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2095_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2095_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2095_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2095_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2095_root_address : std_logic_vector(13 downto 0);
    signal arrayidx82_2074 : std_logic_vector(31 downto 0);
    signal arrayidx87_2097 : std_logic_vector(31 downto 0);
    signal call11_1873 : std_logic_vector(15 downto 0);
    signal call13_1876 : std_logic_vector(15 downto 0);
    signal call14_1879 : std_logic_vector(15 downto 0);
    signal call15_1882 : std_logic_vector(15 downto 0);
    signal call16_1895 : std_logic_vector(15 downto 0);
    signal call18_1907 : std_logic_vector(15 downto 0);
    signal call1_1858 : std_logic_vector(15 downto 0);
    signal call20_1910 : std_logic_vector(15 downto 0);
    signal call22_1913 : std_logic_vector(15 downto 0);
    signal call3_1861 : std_logic_vector(15 downto 0);
    signal call5_1864 : std_logic_vector(15 downto 0);
    signal call7_1867 : std_logic_vector(15 downto 0);
    signal call9_1870 : std_logic_vector(15 downto 0);
    signal call_1855 : std_logic_vector(15 downto 0);
    signal cmp106_2142 : std_logic_vector(0 downto 0);
    signal cmp117_2167 : std_logic_vector(0 downto 0);
    signal cmp_2116 : std_logic_vector(0 downto 0);
    signal conv112_2162 : std_logic_vector(31 downto 0);
    signal conv115_1958 : std_logic_vector(31 downto 0);
    signal conv17_1899 : std_logic_vector(31 downto 0);
    signal conv65_2029 : std_logic_vector(63 downto 0);
    signal conv68_1946 : std_logic_vector(63 downto 0);
    signal conv70_2033 : std_logic_vector(63 downto 0);
    signal conv73_1950 : std_logic_vector(63 downto 0);
    signal conv75_2037 : std_logic_vector(63 downto 0);
    signal conv90_2105 : std_logic_vector(31 downto 0);
    signal conv94_1954 : std_logic_vector(31 downto 0);
    signal conv_1886 : std_logic_vector(31 downto 0);
    signal idxprom86_2090 : std_logic_vector(63 downto 0);
    signal idxprom_2067 : std_logic_vector(63 downto 0);
    signal inc110_2146 : std_logic_vector(15 downto 0);
    signal inc110x_xinput_dim0x_x2_2151 : std_logic_vector(15 downto 0);
    signal inc_2137 : std_logic_vector(15 downto 0);
    signal indvar_1967 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_2200 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_2188 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_1988 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_2182 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_1981 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2158 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_2175 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1974 : std_logic_vector(15 downto 0);
    signal mul54_2020 : std_logic_vector(15 downto 0);
    signal mul76_2042 : std_logic_vector(63 downto 0);
    signal mul78_2052 : std_logic_vector(63 downto 0);
    signal mul_2010 : std_logic_vector(15 downto 0);
    signal ptr_deref_2077_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2077_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2077_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2077_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2077_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2099_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2099_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2099_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2099_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2099_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2099_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_1892 : std_logic_vector(31 downto 0);
    signal shr116132_1964 : std_logic_vector(31 downto 0);
    signal shr131_1920 : std_logic_vector(15 downto 0);
    signal shr81_2063 : std_logic_vector(31 downto 0);
    signal shr85_2084 : std_logic_vector(63 downto 0);
    signal sub48_2015 : std_logic_vector(15 downto 0);
    signal sub61_1942 : std_logic_vector(15 downto 0);
    signal sub62_2025 : std_logic_vector(15 downto 0);
    signal sub_1931 : std_logic_vector(15 downto 0);
    signal tmp1_2000 : std_logic_vector(31 downto 0);
    signal tmp83_2078 : std_logic_vector(63 downto 0);
    signal type_cast_1890_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1918_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1924_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1935_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1962_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1971_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1973_wire : std_logic_vector(31 downto 0);
    signal type_cast_1978_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1980_wire : std_logic_vector(15 downto 0);
    signal type_cast_1985_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1987_wire : std_logic_vector(15 downto 0);
    signal type_cast_1991_wire : std_logic_vector(15 downto 0);
    signal type_cast_1993_wire : std_logic_vector(15 downto 0);
    signal type_cast_1998_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2061_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2082_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2088_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2109_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2127_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2135_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2155_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2178_wire : std_logic_vector(15 downto 0);
    signal type_cast_2181_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2185_wire : std_logic_vector(15 downto 0);
    signal type_cast_2187_wire : std_logic_vector(15 downto 0);
    signal type_cast_2191_wire : std_logic_vector(15 downto 0);
    signal type_cast_2193_wire : std_logic_vector(15 downto 0);
    signal type_cast_2198_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2206_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_2072_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2072_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2072_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2072_resized_base_address <= "00000000000000";
    array_obj_ref_2095_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2095_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2095_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2095_resized_base_address <= "00000000000000";
    ptr_deref_2077_word_offset_0 <= "00000000000000";
    ptr_deref_2099_word_offset_0 <= "00000000000000";
    type_cast_1890_wire_constant <= "00000000000000000000000000010000";
    type_cast_1918_wire_constant <= "0000000000000010";
    type_cast_1924_wire_constant <= "1111111111111111";
    type_cast_1935_wire_constant <= "1111111111111111";
    type_cast_1962_wire_constant <= "00000000000000000000000000000001";
    type_cast_1971_wire_constant <= "00000000000000000000000000000000";
    type_cast_1978_wire_constant <= "0000000000000000";
    type_cast_1985_wire_constant <= "0000000000000000";
    type_cast_1998_wire_constant <= "00000000000000000000000000000100";
    type_cast_2061_wire_constant <= "00000000000000000000000000000010";
    type_cast_2082_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_2088_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_2109_wire_constant <= "00000000000000000000000000000100";
    type_cast_2127_wire_constant <= "0000000000000100";
    type_cast_2135_wire_constant <= "0000000000000001";
    type_cast_2155_wire_constant <= "0000000000000000";
    type_cast_2181_wire_constant <= "0000000000000000";
    type_cast_2198_wire_constant <= "00000000000000000000000000000001";
    type_cast_2206_wire_constant <= "0000000000000001";
    phi_stmt_1967: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1971_wire_constant & type_cast_1973_wire;
      req <= phi_stmt_1967_req_0 & phi_stmt_1967_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1967",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1967_ack_0,
          idata => idata,
          odata => indvar_1967,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1967
    phi_stmt_1974: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1978_wire_constant & type_cast_1980_wire;
      req <= phi_stmt_1974_req_0 & phi_stmt_1974_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1974",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1974_ack_0,
          idata => idata,
          odata => input_dim2x_x1_1974,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1974
    phi_stmt_1981: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1985_wire_constant & type_cast_1987_wire;
      req <= phi_stmt_1981_req_0 & phi_stmt_1981_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1981",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1981_ack_0,
          idata => idata,
          odata => input_dim1x_x1_1981,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1981
    phi_stmt_1988: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1991_wire & type_cast_1993_wire;
      req <= phi_stmt_1988_req_0 & phi_stmt_1988_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1988",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1988_ack_0,
          idata => idata,
          odata => input_dim0x_x2_1988,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1988
    phi_stmt_2175: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2178_wire & type_cast_2181_wire_constant;
      req <= phi_stmt_2175_req_0 & phi_stmt_2175_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2175",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2175_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_2175,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2175
    phi_stmt_2182: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2185_wire & type_cast_2187_wire;
      req <= phi_stmt_2182_req_0 & phi_stmt_2182_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2182",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2182_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_2182,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2182
    phi_stmt_2188: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2191_wire & type_cast_2193_wire;
      req <= phi_stmt_2188_req_0 & phi_stmt_2188_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2188",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2188_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_2188,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2188
    -- flow-through select operator MUX_2157_inst
    input_dim1x_x2_2158 <= type_cast_2155_wire_constant when (cmp106_2142(0) /=  '0') else inc_2137;
    addr_of_2073_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2073_final_reg_req_0;
      addr_of_2073_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2073_final_reg_req_1;
      addr_of_2073_final_reg_ack_1<= rack(0);
      addr_of_2073_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2073_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2072_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx82_2074,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2096_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2096_final_reg_req_0;
      addr_of_2096_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2096_final_reg_req_1;
      addr_of_2096_final_reg_ack_1<= rack(0);
      addr_of_2096_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2096_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2095_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx87_2097,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1885_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1885_inst_req_0;
      type_cast_1885_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1885_inst_req_1;
      type_cast_1885_inst_ack_1<= rack(0);
      type_cast_1885_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1885_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_1882,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1886,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1898_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1898_inst_req_0;
      type_cast_1898_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1898_inst_req_1;
      type_cast_1898_inst_ack_1<= rack(0);
      type_cast_1898_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1898_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_1895,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_1899,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1945_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1945_inst_req_0;
      type_cast_1945_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1945_inst_req_1;
      type_cast_1945_inst_ack_1<= rack(0);
      type_cast_1945_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1945_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_1913,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv68_1946,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1949_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1949_inst_req_0;
      type_cast_1949_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1949_inst_req_1;
      type_cast_1949_inst_ack_1<= rack(0);
      type_cast_1949_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1949_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_1910,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_1950,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1953_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1953_inst_req_0;
      type_cast_1953_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1953_inst_req_1;
      type_cast_1953_inst_ack_1<= rack(0);
      type_cast_1953_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1953_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_1861,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv94_1954,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1957_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1957_inst_req_0;
      type_cast_1957_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1957_inst_req_1;
      type_cast_1957_inst_ack_1<= rack(0);
      type_cast_1957_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1957_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1855,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv115_1958,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1973_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1973_inst_req_0;
      type_cast_1973_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1973_inst_req_1;
      type_cast_1973_inst_ack_1<= rack(0);
      type_cast_1973_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1973_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2200,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1973_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1980_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1980_inst_req_0;
      type_cast_1980_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1980_inst_req_1;
      type_cast_1980_inst_ack_1<= rack(0);
      type_cast_1980_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1980_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_2175,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1980_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1987_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1987_inst_req_0;
      type_cast_1987_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1987_inst_req_1;
      type_cast_1987_inst_ack_1<= rack(0);
      type_cast_1987_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1987_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_2182,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1987_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1991_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1991_inst_req_0;
      type_cast_1991_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1991_inst_req_1;
      type_cast_1991_inst_ack_1<= rack(0);
      type_cast_1991_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1991_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr131_1920,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1991_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1993_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1993_inst_req_0;
      type_cast_1993_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1993_inst_req_1;
      type_cast_1993_inst_ack_1<= rack(0);
      type_cast_1993_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1993_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_2188,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1993_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2028_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2028_inst_req_0;
      type_cast_2028_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2028_inst_req_1;
      type_cast_2028_inst_ack_1<= rack(0);
      type_cast_2028_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2028_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1974,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_2029,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2032_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2032_inst_req_0;
      type_cast_2032_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2032_inst_req_1;
      type_cast_2032_inst_ack_1<= rack(0);
      type_cast_2032_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2032_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub62_2025,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_2033,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2036_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2036_inst_req_0;
      type_cast_2036_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2036_inst_req_1;
      type_cast_2036_inst_ack_1<= rack(0);
      type_cast_2036_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2036_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub48_2015,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_2037,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2066_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2066_inst_req_0;
      type_cast_2066_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2066_inst_req_1;
      type_cast_2066_inst_ack_1<= rack(0);
      type_cast_2066_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2066_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr81_2063,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2067,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2104_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2104_inst_req_0;
      type_cast_2104_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2104_inst_req_1;
      type_cast_2104_inst_ack_1<= rack(0);
      type_cast_2104_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2104_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1974,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_2105,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2145_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2145_inst_req_0;
      type_cast_2145_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2145_inst_req_1;
      type_cast_2145_inst_ack_1<= rack(0);
      type_cast_2145_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2145_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp106_2142,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc110_2146,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2161_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2161_inst_req_0;
      type_cast_2161_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2161_inst_req_1;
      type_cast_2161_inst_ack_1<= rack(0);
      type_cast_2161_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2161_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc110x_xinput_dim0x_x2_2151,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv112_2162,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2178_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2178_inst_req_0;
      type_cast_2178_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2178_inst_req_1;
      type_cast_2178_inst_ack_1<= rack(0);
      type_cast_2178_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2178_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add98_2129,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2178_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2185_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2185_inst_req_0;
      type_cast_2185_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2185_inst_req_1;
      type_cast_2185_inst_ack_1<= rack(0);
      type_cast_2185_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2185_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2158,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2185_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2187_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2187_inst_req_0;
      type_cast_2187_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2187_inst_req_1;
      type_cast_2187_inst_ack_1<= rack(0);
      type_cast_2187_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2187_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_1981,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2187_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2191_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2191_inst_req_0;
      type_cast_2191_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2191_inst_req_1;
      type_cast_2191_inst_ack_1<= rack(0);
      type_cast_2191_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2191_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_1988,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2191_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2193_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2193_inst_req_0;
      type_cast_2193_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2193_inst_req_1;
      type_cast_2193_inst_ack_1<= rack(0);
      type_cast_2193_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2193_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc110x_xinput_dim0x_x2_2151,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2193_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_2072_index_1_rename
    process(R_idxprom_2071_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2071_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2071_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2072_index_1_resize
    process(idxprom_2067) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2067;
      ov := iv(13 downto 0);
      R_idxprom_2071_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2072_root_address_inst
    process(array_obj_ref_2072_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2072_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2072_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2095_index_1_rename
    process(R_idxprom86_2094_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom86_2094_resized;
      ov(13 downto 0) := iv;
      R_idxprom86_2094_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2095_index_1_resize
    process(idxprom86_2090) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom86_2090;
      ov := iv(13 downto 0);
      R_idxprom86_2094_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2095_root_address_inst
    process(array_obj_ref_2095_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2095_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2095_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2077_addr_0
    process(ptr_deref_2077_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2077_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2077_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2077_base_resize
    process(arrayidx82_2074) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx82_2074;
      ov := iv(13 downto 0);
      ptr_deref_2077_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2077_gather_scatter
    process(ptr_deref_2077_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2077_data_0;
      ov(63 downto 0) := iv;
      tmp83_2078 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2077_root_address_inst
    process(ptr_deref_2077_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2077_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2077_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2099_addr_0
    process(ptr_deref_2099_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2099_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2099_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2099_base_resize
    process(arrayidx87_2097) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx87_2097;
      ov := iv(13 downto 0);
      ptr_deref_2099_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2099_gather_scatter
    process(tmp83_2078) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp83_2078;
      ov(63 downto 0) := iv;
      ptr_deref_2099_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2099_root_address_inst
    process(ptr_deref_2099_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2099_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2099_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2117_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2116;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2117_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2117_branch_req_0,
          ack0 => if_stmt_2117_branch_ack_0,
          ack1 => if_stmt_2117_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2168_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp117_2167;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2168_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2168_branch_req_0,
          ack0 => if_stmt_2168_branch_ack_0,
          ack1 => if_stmt_2168_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1925_inst
    process(call7_1867) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_1867, type_cast_1924_wire_constant, tmp_var);
      add45_1926 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1936_inst
    process(call9_1870) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_1870, type_cast_1935_wire_constant, tmp_var);
      add58_1937 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2014_inst
    process(sub_1931, mul_2010) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_1931, mul_2010, tmp_var);
      sub48_2015 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2024_inst
    process(sub61_1942, mul54_2020) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub61_1942, mul54_2020, tmp_var);
      sub62_2025 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2128_inst
    process(input_dim2x_x1_1974) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_1974, type_cast_2127_wire_constant, tmp_var);
      add98_2129 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2136_inst
    process(input_dim1x_x1_1981) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_1981, type_cast_2135_wire_constant, tmp_var);
      inc_2137 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2150_inst
    process(inc110_2146, input_dim0x_x2_1988) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc110_2146, input_dim0x_x2_1988, tmp_var);
      inc110x_xinput_dim0x_x2_2151 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2004_inst
    process(add_1904, tmp1_2000) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_1904, tmp1_2000, tmp_var);
      add_src_0x_x0_2005 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2110_inst
    process(conv90_2105) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv90_2105, type_cast_2109_wire_constant, tmp_var);
      add91_2111 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2199_inst
    process(indvar_1967) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1967, type_cast_2198_wire_constant, tmp_var);
      indvarx_xnext_2200 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2046_inst
    process(mul76_2042, conv70_2033) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul76_2042, conv70_2033, tmp_var);
      add77_2047 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2056_inst
    process(mul78_2052, conv65_2029) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul78_2052, conv65_2029, tmp_var);
      add79_2057 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2089_inst
    process(shr85_2084) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr85_2084, type_cast_2088_wire_constant, tmp_var);
      idxprom86_2090 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2141_inst
    process(inc_2137, call1_1858) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_2137, call1_1858, tmp_var);
      cmp106_2142 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2166_inst
    process(conv112_2162, shr116132_1964) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv112_2162, shr116132_1964, tmp_var);
      cmp117_2167 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_1919_inst
    process(call_1855) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_1855, type_cast_1918_wire_constant, tmp_var);
      shr131_1920 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1963_inst
    process(conv115_1958) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv115_1958, type_cast_1962_wire_constant, tmp_var);
      shr116132_1964 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2062_inst
    process(add_src_0x_x0_2005) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_2005, type_cast_2061_wire_constant, tmp_var);
      shr81_2063 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2083_inst
    process(add79_2057) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add79_2057, type_cast_2082_wire_constant, tmp_var);
      shr85_2084 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2009_inst
    process(input_dim0x_x2_1988, call13_1876) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x2_1988, call13_1876, tmp_var);
      mul_2010 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2019_inst
    process(input_dim1x_x1_1981, call13_1876) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_1981, call13_1876, tmp_var);
      mul54_2020 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1999_inst
    process(indvar_1967) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_1967, type_cast_1998_wire_constant, tmp_var);
      tmp1_2000 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2041_inst
    process(conv75_2037, conv73_1950) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv75_2037, conv73_1950, tmp_var);
      mul76_2042 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2051_inst
    process(add77_2047, conv68_1946) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add77_2047, conv68_1946, tmp_var);
      mul78_2052 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1903_inst
    process(shl_1892, conv17_1899) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_1892, conv17_1899, tmp_var);
      add_1904 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1891_inst
    process(conv_1886) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_1886, type_cast_1890_wire_constant, tmp_var);
      shl_1892 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1930_inst
    process(add45_1926, call14_1879) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add45_1926, call14_1879, tmp_var);
      sub_1931 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1941_inst
    process(add58_1937, call14_1879) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add58_1937, call14_1879, tmp_var);
      sub61_1942 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2115_inst
    process(add91_2111, conv94_1954) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add91_2111, conv94_1954, tmp_var);
      cmp_2116 <= tmp_var; --
    end process;
    -- shared split operator group (29) : array_obj_ref_2072_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2071_scaled;
      array_obj_ref_2072_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2072_index_offset_req_0;
      array_obj_ref_2072_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2072_index_offset_req_1;
      array_obj_ref_2072_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : array_obj_ref_2095_index_offset 
    ApIntAdd_group_30: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom86_2094_scaled;
      array_obj_ref_2095_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2095_index_offset_req_0;
      array_obj_ref_2095_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2095_index_offset_req_1;
      array_obj_ref_2095_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_30_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_30_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_30",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared load operator group (0) : ptr_deref_2077_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2077_load_0_req_0;
      ptr_deref_2077_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2077_load_0_req_1;
      ptr_deref_2077_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2077_word_address_0;
      ptr_deref_2077_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_2099_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2099_store_0_req_0;
      ptr_deref_2099_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2099_store_0_req_1;
      ptr_deref_2099_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2099_word_address_0;
      data_in <= ptr_deref_2099_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block1_start_1912_inst RPIPE_Block1_start_1909_inst RPIPE_Block1_start_1906_inst RPIPE_Block1_start_1894_inst RPIPE_Block1_start_1881_inst RPIPE_Block1_start_1878_inst RPIPE_Block1_start_1875_inst RPIPE_Block1_start_1872_inst RPIPE_Block1_start_1869_inst RPIPE_Block1_start_1866_inst RPIPE_Block1_start_1863_inst RPIPE_Block1_start_1860_inst RPIPE_Block1_start_1857_inst RPIPE_Block1_start_1854_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block1_start_1912_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block1_start_1909_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block1_start_1906_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block1_start_1894_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block1_start_1881_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block1_start_1878_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block1_start_1875_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block1_start_1872_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block1_start_1869_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block1_start_1866_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block1_start_1863_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block1_start_1860_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block1_start_1857_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block1_start_1854_inst_req_0;
      RPIPE_Block1_start_1912_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block1_start_1909_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block1_start_1906_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block1_start_1894_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block1_start_1881_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block1_start_1878_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block1_start_1875_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block1_start_1872_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block1_start_1869_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block1_start_1866_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block1_start_1863_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block1_start_1860_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block1_start_1857_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block1_start_1854_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block1_start_1912_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block1_start_1909_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block1_start_1906_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block1_start_1894_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block1_start_1881_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block1_start_1878_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block1_start_1875_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block1_start_1872_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block1_start_1869_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block1_start_1866_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block1_start_1863_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block1_start_1860_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block1_start_1857_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block1_start_1854_inst_req_1;
      RPIPE_Block1_start_1912_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block1_start_1909_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block1_start_1906_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block1_start_1894_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block1_start_1881_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block1_start_1878_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block1_start_1875_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block1_start_1872_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block1_start_1869_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block1_start_1866_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block1_start_1863_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block1_start_1860_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block1_start_1857_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block1_start_1854_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call22_1913 <= data_out(223 downto 208);
      call20_1910 <= data_out(207 downto 192);
      call18_1907 <= data_out(191 downto 176);
      call16_1895 <= data_out(175 downto 160);
      call15_1882 <= data_out(159 downto 144);
      call14_1879 <= data_out(143 downto 128);
      call13_1876 <= data_out(127 downto 112);
      call11_1873 <= data_out(111 downto 96);
      call9_1870 <= data_out(95 downto 80);
      call7_1867 <= data_out(79 downto 64);
      call5_1864 <= data_out(63 downto 48);
      call3_1861 <= data_out(47 downto 32);
      call1_1858 <= data_out(31 downto 16);
      call_1855 <= data_out(15 downto 0);
      Block1_start_read_0_gI: SplitGuardInterface generic map(name => "Block1_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_start_read_0: InputPortRevised -- 
        generic map ( name => "Block1_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_start_pipe_read_req(0),
          oack => Block1_start_pipe_read_ack(0),
          odata => Block1_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block1_done_2204_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block1_done_2204_inst_req_0;
      WPIPE_Block1_done_2204_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block1_done_2204_inst_req_1;
      WPIPE_Block1_done_2204_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2206_wire_constant;
      Block1_done_write_0_gI: SplitGuardInterface generic map(name => "Block1_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block1_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_done_pipe_write_req(0),
          oack => Block1_done_pipe_write_ack(0),
          odata => Block1_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeB_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeC is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeC;
architecture convTransposeC_arch of convTransposeC is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeC_CP_5782_start: Boolean;
  signal convTransposeC_CP_5782_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block2_start_2233_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2221_inst_ack_1 : boolean;
  signal type_cast_2259_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2221_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2224_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2239_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2233_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2239_inst_req_0 : boolean;
  signal type_cast_2246_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2233_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2255_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2267_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2227_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2270_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2255_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2230_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2273_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2273_inst_req_0 : boolean;
  signal type_cast_2246_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2230_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2227_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2227_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2227_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2239_inst_req_1 : boolean;
  signal type_cast_2259_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2236_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2239_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2236_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2236_inst_ack_0 : boolean;
  signal type_cast_2246_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2221_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2242_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2255_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2255_inst_ack_1 : boolean;
  signal type_cast_2246_inst_ack_0 : boolean;
  signal type_cast_2259_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2267_inst_req_0 : boolean;
  signal type_cast_2306_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2242_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2242_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2233_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2230_inst_ack_0 : boolean;
  signal type_cast_2259_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2242_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2267_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2224_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2230_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2224_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2267_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2236_inst_req_1 : boolean;
  signal type_cast_2306_inst_req_1 : boolean;
  signal type_cast_2306_inst_ack_1 : boolean;
  signal type_cast_2314_inst_req_1 : boolean;
  signal type_cast_2314_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2270_inst_req_1 : boolean;
  signal type_cast_2310_inst_req_1 : boolean;
  signal type_cast_2310_inst_ack_1 : boolean;
  signal type_cast_2310_inst_req_0 : boolean;
  signal type_cast_2310_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2273_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2270_inst_ack_0 : boolean;
  signal type_cast_2314_inst_req_0 : boolean;
  signal type_cast_2314_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2273_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2270_inst_req_0 : boolean;
  signal type_cast_2306_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2224_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2221_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2215_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2215_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2215_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2215_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2218_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2218_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2218_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2218_inst_ack_1 : boolean;
  signal type_cast_2318_inst_req_0 : boolean;
  signal type_cast_2318_inst_ack_0 : boolean;
  signal type_cast_2318_inst_req_1 : boolean;
  signal type_cast_2318_inst_ack_1 : boolean;
  signal type_cast_2400_inst_req_0 : boolean;
  signal type_cast_2400_inst_ack_0 : boolean;
  signal type_cast_2400_inst_req_1 : boolean;
  signal type_cast_2400_inst_ack_1 : boolean;
  signal type_cast_2404_inst_req_0 : boolean;
  signal type_cast_2404_inst_ack_0 : boolean;
  signal type_cast_2404_inst_req_1 : boolean;
  signal type_cast_2404_inst_ack_1 : boolean;
  signal type_cast_2408_inst_req_0 : boolean;
  signal type_cast_2408_inst_ack_0 : boolean;
  signal type_cast_2408_inst_req_1 : boolean;
  signal type_cast_2408_inst_ack_1 : boolean;
  signal type_cast_2438_inst_req_0 : boolean;
  signal type_cast_2438_inst_ack_0 : boolean;
  signal type_cast_2438_inst_req_1 : boolean;
  signal type_cast_2438_inst_ack_1 : boolean;
  signal array_obj_ref_2444_index_offset_req_0 : boolean;
  signal array_obj_ref_2444_index_offset_ack_0 : boolean;
  signal array_obj_ref_2444_index_offset_req_1 : boolean;
  signal array_obj_ref_2444_index_offset_ack_1 : boolean;
  signal addr_of_2445_final_reg_req_0 : boolean;
  signal addr_of_2445_final_reg_ack_0 : boolean;
  signal addr_of_2445_final_reg_req_1 : boolean;
  signal addr_of_2445_final_reg_ack_1 : boolean;
  signal ptr_deref_2449_load_0_req_0 : boolean;
  signal ptr_deref_2449_load_0_ack_0 : boolean;
  signal ptr_deref_2449_load_0_req_1 : boolean;
  signal ptr_deref_2449_load_0_ack_1 : boolean;
  signal array_obj_ref_2467_index_offset_req_0 : boolean;
  signal array_obj_ref_2467_index_offset_ack_0 : boolean;
  signal array_obj_ref_2467_index_offset_req_1 : boolean;
  signal array_obj_ref_2467_index_offset_ack_1 : boolean;
  signal addr_of_2468_final_reg_req_0 : boolean;
  signal addr_of_2468_final_reg_ack_0 : boolean;
  signal addr_of_2468_final_reg_req_1 : boolean;
  signal addr_of_2468_final_reg_ack_1 : boolean;
  signal ptr_deref_2471_store_0_req_0 : boolean;
  signal ptr_deref_2471_store_0_ack_0 : boolean;
  signal ptr_deref_2471_store_0_req_1 : boolean;
  signal ptr_deref_2471_store_0_ack_1 : boolean;
  signal type_cast_2476_inst_req_0 : boolean;
  signal type_cast_2476_inst_ack_0 : boolean;
  signal type_cast_2476_inst_req_1 : boolean;
  signal type_cast_2476_inst_ack_1 : boolean;
  signal if_stmt_2489_branch_req_0 : boolean;
  signal if_stmt_2489_branch_ack_1 : boolean;
  signal if_stmt_2489_branch_ack_0 : boolean;
  signal type_cast_2517_inst_req_0 : boolean;
  signal type_cast_2517_inst_ack_0 : boolean;
  signal type_cast_2517_inst_req_1 : boolean;
  signal type_cast_2517_inst_ack_1 : boolean;
  signal type_cast_2533_inst_req_0 : boolean;
  signal type_cast_2533_inst_ack_0 : boolean;
  signal type_cast_2533_inst_req_1 : boolean;
  signal type_cast_2533_inst_ack_1 : boolean;
  signal if_stmt_2540_branch_req_0 : boolean;
  signal if_stmt_2540_branch_ack_1 : boolean;
  signal if_stmt_2540_branch_ack_0 : boolean;
  signal WPIPE_Block2_done_2576_inst_req_0 : boolean;
  signal WPIPE_Block2_done_2576_inst_ack_0 : boolean;
  signal WPIPE_Block2_done_2576_inst_req_1 : boolean;
  signal WPIPE_Block2_done_2576_inst_ack_1 : boolean;
  signal phi_stmt_2339_req_0 : boolean;
  signal phi_stmt_2346_req_0 : boolean;
  signal phi_stmt_2353_req_1 : boolean;
  signal type_cast_2365_inst_req_0 : boolean;
  signal type_cast_2365_inst_ack_0 : boolean;
  signal type_cast_2365_inst_req_1 : boolean;
  signal type_cast_2365_inst_ack_1 : boolean;
  signal phi_stmt_2360_req_1 : boolean;
  signal type_cast_2345_inst_req_0 : boolean;
  signal type_cast_2345_inst_ack_0 : boolean;
  signal type_cast_2345_inst_req_1 : boolean;
  signal type_cast_2345_inst_ack_1 : boolean;
  signal phi_stmt_2339_req_1 : boolean;
  signal type_cast_2352_inst_req_0 : boolean;
  signal type_cast_2352_inst_ack_0 : boolean;
  signal type_cast_2352_inst_req_1 : boolean;
  signal type_cast_2352_inst_ack_1 : boolean;
  signal phi_stmt_2346_req_1 : boolean;
  signal type_cast_2356_inst_req_0 : boolean;
  signal type_cast_2356_inst_ack_0 : boolean;
  signal type_cast_2356_inst_req_1 : boolean;
  signal type_cast_2356_inst_ack_1 : boolean;
  signal phi_stmt_2353_req_0 : boolean;
  signal type_cast_2363_inst_req_0 : boolean;
  signal type_cast_2363_inst_ack_0 : boolean;
  signal type_cast_2363_inst_req_1 : boolean;
  signal type_cast_2363_inst_ack_1 : boolean;
  signal phi_stmt_2360_req_0 : boolean;
  signal phi_stmt_2339_ack_0 : boolean;
  signal phi_stmt_2346_ack_0 : boolean;
  signal phi_stmt_2353_ack_0 : boolean;
  signal phi_stmt_2360_ack_0 : boolean;
  signal phi_stmt_2547_req_1 : boolean;
  signal type_cast_2557_inst_req_0 : boolean;
  signal type_cast_2557_inst_ack_0 : boolean;
  signal type_cast_2557_inst_req_1 : boolean;
  signal type_cast_2557_inst_ack_1 : boolean;
  signal phi_stmt_2554_req_0 : boolean;
  signal type_cast_2563_inst_req_0 : boolean;
  signal type_cast_2563_inst_ack_0 : boolean;
  signal type_cast_2563_inst_req_1 : boolean;
  signal type_cast_2563_inst_ack_1 : boolean;
  signal phi_stmt_2560_req_0 : boolean;
  signal type_cast_2550_inst_req_0 : boolean;
  signal type_cast_2550_inst_ack_0 : boolean;
  signal type_cast_2550_inst_req_1 : boolean;
  signal type_cast_2550_inst_ack_1 : boolean;
  signal phi_stmt_2547_req_0 : boolean;
  signal type_cast_2559_inst_req_0 : boolean;
  signal type_cast_2559_inst_ack_0 : boolean;
  signal type_cast_2559_inst_req_1 : boolean;
  signal type_cast_2559_inst_ack_1 : boolean;
  signal phi_stmt_2554_req_1 : boolean;
  signal type_cast_2565_inst_req_0 : boolean;
  signal type_cast_2565_inst_ack_0 : boolean;
  signal type_cast_2565_inst_req_1 : boolean;
  signal type_cast_2565_inst_ack_1 : boolean;
  signal phi_stmt_2560_req_1 : boolean;
  signal phi_stmt_2547_ack_0 : boolean;
  signal phi_stmt_2554_ack_0 : boolean;
  signal phi_stmt_2560_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeC_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeC_CP_5782_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeC_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_5782_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeC_CP_5782_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_5782_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeC_CP_5782: Block -- control-path 
    signal convTransposeC_CP_5782_elements: BooleanArray(127 downto 0);
    -- 
  begin -- 
    convTransposeC_CP_5782_elements(0) <= convTransposeC_CP_5782_start;
    convTransposeC_CP_5782_symbol <= convTransposeC_CP_5782_elements(78);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/type_cast_2246_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/type_cast_2259_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/type_cast_2246_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/type_cast_2259_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/type_cast_2259_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/type_cast_2246_update_start_
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2213/$entry
      -- CP-element group 0: 	 branch_block_stmt_2213/branch_block_stmt_2213__entry__
      -- CP-element group 0: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274__entry__
      -- CP-element group 0: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/$entry
      -- CP-element group 0: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2215_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2215_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2215_Sample/rr
      -- 
    cr_5975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(0), ack => type_cast_2246_inst_req_1); -- 
    cr_6003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(0), ack => type_cast_2259_inst_req_1); -- 
    rr_5830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(0), ack => RPIPE_Block2_start_2215_inst_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	127 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	86 
    -- CP-element group 1: 	87 
    -- CP-element group 1: 	89 
    -- CP-element group 1: 	90 
    -- CP-element group 1: 	92 
    -- CP-element group 1: 	93 
    -- CP-element group 1: 	95 
    -- CP-element group 1: 	96 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_2213/merge_stmt_2546__exit__
      -- CP-element group 1: 	 branch_block_stmt_2213/assign_stmt_2572__entry__
      -- CP-element group 1: 	 branch_block_stmt_2213/assign_stmt_2572__exit__
      -- CP-element group 1: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_2213/assign_stmt_2572/$entry
      -- CP-element group 1: 	 branch_block_stmt_2213/assign_stmt_2572/$exit
      -- CP-element group 1: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2339/$entry
      -- CP-element group 1: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2339/phi_stmt_2339_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2339/phi_stmt_2339_sources/type_cast_2345/$entry
      -- CP-element group 1: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2339/phi_stmt_2339_sources/type_cast_2345/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2339/phi_stmt_2339_sources/type_cast_2345/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2339/phi_stmt_2339_sources/type_cast_2345/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2339/phi_stmt_2339_sources/type_cast_2345/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2339/phi_stmt_2339_sources/type_cast_2345/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2346/$entry
      -- CP-element group 1: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2346/phi_stmt_2346_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2346/phi_stmt_2346_sources/type_cast_2352/$entry
      -- CP-element group 1: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2346/phi_stmt_2346_sources/type_cast_2352/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2346/phi_stmt_2346_sources/type_cast_2352/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2346/phi_stmt_2346_sources/type_cast_2352/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2346/phi_stmt_2346_sources/type_cast_2352/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2346/phi_stmt_2346_sources/type_cast_2352/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2353/$entry
      -- CP-element group 1: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2353/phi_stmt_2353_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2353/phi_stmt_2353_sources/type_cast_2356/$entry
      -- CP-element group 1: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2353/phi_stmt_2353_sources/type_cast_2356/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2353/phi_stmt_2353_sources/type_cast_2356/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2353/phi_stmt_2353_sources/type_cast_2356/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2353/phi_stmt_2353_sources/type_cast_2356/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2353/phi_stmt_2353_sources/type_cast_2356/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2360/$entry
      -- CP-element group 1: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2360/phi_stmt_2360_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2360/phi_stmt_2360_sources/type_cast_2363/$entry
      -- CP-element group 1: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2360/phi_stmt_2360_sources/type_cast_2363/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2360/phi_stmt_2360_sources/type_cast_2363/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2360/phi_stmt_2360_sources/type_cast_2363/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2360/phi_stmt_2360_sources/type_cast_2363/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2360/phi_stmt_2360_sources/type_cast_2363/SplitProtocol/Update/cr
      -- 
    rr_6531_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6531_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(1), ack => type_cast_2345_inst_req_0); -- 
    cr_6536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(1), ack => type_cast_2345_inst_req_1); -- 
    rr_6554_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6554_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(1), ack => type_cast_2352_inst_req_0); -- 
    cr_6559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(1), ack => type_cast_2352_inst_req_1); -- 
    rr_6577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(1), ack => type_cast_2356_inst_req_0); -- 
    cr_6582_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6582_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(1), ack => type_cast_2356_inst_req_1); -- 
    rr_6600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(1), ack => type_cast_2363_inst_req_0); -- 
    cr_6605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(1), ack => type_cast_2363_inst_req_1); -- 
    convTransposeC_CP_5782_elements(1) <= convTransposeC_CP_5782_elements(127);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2215_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2215_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2215_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2215_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2215_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2215_Update/cr
      -- 
    ra_5831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2215_inst_ack_0, ack => convTransposeC_CP_5782_elements(2)); -- 
    cr_5835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(2), ack => RPIPE_Block2_start_2215_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2215_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2215_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2215_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2218_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2218_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2218_Sample/rr
      -- 
    ca_5836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2215_inst_ack_1, ack => convTransposeC_CP_5782_elements(3)); -- 
    rr_5844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(3), ack => RPIPE_Block2_start_2218_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2218_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2218_update_start_
      -- CP-element group 4: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2218_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2218_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2218_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2218_Update/cr
      -- 
    ra_5845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2218_inst_ack_0, ack => convTransposeC_CP_5782_elements(4)); -- 
    cr_5849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(4), ack => RPIPE_Block2_start_2218_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2221_Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2221_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2218_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2218_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2218_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2221_sample_start_
      -- 
    ca_5850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2218_inst_ack_1, ack => convTransposeC_CP_5782_elements(5)); -- 
    rr_5858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(5), ack => RPIPE_Block2_start_2221_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2221_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2221_Update/cr
      -- CP-element group 6: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2221_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2221_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2221_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2221_update_start_
      -- 
    ra_5859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2221_inst_ack_0, ack => convTransposeC_CP_5782_elements(6)); -- 
    cr_5863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(6), ack => RPIPE_Block2_start_2221_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2221_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2221_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2224_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2224_Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2224_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2221_update_completed_
      -- 
    ca_5864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2221_inst_ack_1, ack => convTransposeC_CP_5782_elements(7)); -- 
    rr_5872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(7), ack => RPIPE_Block2_start_2224_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2224_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2224_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2224_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2224_update_start_
      -- CP-element group 8: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2224_Update/cr
      -- CP-element group 8: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2224_Sample/$exit
      -- 
    ra_5873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2224_inst_ack_0, ack => convTransposeC_CP_5782_elements(8)); -- 
    cr_5877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(8), ack => RPIPE_Block2_start_2224_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2227_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2227_Sample/rr
      -- CP-element group 9: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2224_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2224_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2224_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2227_sample_start_
      -- 
    ca_5878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2224_inst_ack_1, ack => convTransposeC_CP_5782_elements(9)); -- 
    rr_5886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(9), ack => RPIPE_Block2_start_2227_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2227_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2227_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2227_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2227_update_start_
      -- CP-element group 10: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2227_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2227_sample_completed_
      -- 
    ra_5887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2227_inst_ack_0, ack => convTransposeC_CP_5782_elements(10)); -- 
    cr_5891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(10), ack => RPIPE_Block2_start_2227_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2227_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2230_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2227_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2230_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2230_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2227_Update/ca
      -- 
    ca_5892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2227_inst_ack_1, ack => convTransposeC_CP_5782_elements(11)); -- 
    rr_5900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(11), ack => RPIPE_Block2_start_2230_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2230_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2230_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2230_Update/cr
      -- CP-element group 12: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2230_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2230_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2230_update_start_
      -- 
    ra_5901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2230_inst_ack_0, ack => convTransposeC_CP_5782_elements(12)); -- 
    cr_5905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(12), ack => RPIPE_Block2_start_2230_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2233_Sample/rr
      -- CP-element group 13: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2230_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2230_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2230_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2233_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2233_sample_start_
      -- 
    ca_5906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2230_inst_ack_1, ack => convTransposeC_CP_5782_elements(13)); -- 
    rr_5914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(13), ack => RPIPE_Block2_start_2233_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2233_Update/cr
      -- CP-element group 14: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2233_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2233_update_start_
      -- CP-element group 14: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2233_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2233_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2233_Sample/$exit
      -- 
    ra_5915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2233_inst_ack_0, ack => convTransposeC_CP_5782_elements(14)); -- 
    cr_5919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(14), ack => RPIPE_Block2_start_2233_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2233_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2236_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2233_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2236_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2233_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2236_Sample/$entry
      -- 
    ca_5920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2233_inst_ack_1, ack => convTransposeC_CP_5782_elements(15)); -- 
    rr_5928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(15), ack => RPIPE_Block2_start_2236_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2236_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2236_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2236_update_start_
      -- CP-element group 16: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2236_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2236_Update/cr
      -- CP-element group 16: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2236_Update/$entry
      -- 
    ra_5929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2236_inst_ack_0, ack => convTransposeC_CP_5782_elements(16)); -- 
    cr_5933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(16), ack => RPIPE_Block2_start_2236_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2239_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2239_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2239_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2236_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2236_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2236_update_completed_
      -- 
    ca_5934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2236_inst_ack_1, ack => convTransposeC_CP_5782_elements(17)); -- 
    rr_5942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(17), ack => RPIPE_Block2_start_2239_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2239_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2239_update_start_
      -- CP-element group 18: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2239_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2239_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2239_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2239_Update/cr
      -- 
    ra_5943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2239_inst_ack_0, ack => convTransposeC_CP_5782_elements(18)); -- 
    cr_5947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(18), ack => RPIPE_Block2_start_2239_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2239_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2239_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2239_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2242_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2242_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2242_Sample/rr
      -- 
    ca_5948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2239_inst_ack_1, ack => convTransposeC_CP_5782_elements(19)); -- 
    rr_5956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(19), ack => RPIPE_Block2_start_2242_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2242_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2242_update_start_
      -- CP-element group 20: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2242_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2242_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2242_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2242_Update/cr
      -- 
    ra_5957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2242_inst_ack_0, ack => convTransposeC_CP_5782_elements(20)); -- 
    cr_5961_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5961_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(20), ack => RPIPE_Block2_start_2242_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/type_cast_2246_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2255_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2255_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2255_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2242_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/type_cast_2246_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2242_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2242_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/type_cast_2246_sample_start_
      -- 
    ca_5962_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2242_inst_ack_1, ack => convTransposeC_CP_5782_elements(21)); -- 
    rr_5970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(21), ack => type_cast_2246_inst_req_0); -- 
    rr_5984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(21), ack => RPIPE_Block2_start_2255_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/type_cast_2246_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/type_cast_2246_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/type_cast_2246_sample_completed_
      -- 
    ra_5971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2246_inst_ack_0, ack => convTransposeC_CP_5782_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/type_cast_2246_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/type_cast_2246_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/type_cast_2246_Update/ca
      -- 
    ca_5976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2246_inst_ack_1, ack => convTransposeC_CP_5782_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2255_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2255_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2255_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2255_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2255_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2255_update_start_
      -- 
    ra_5985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2255_inst_ack_0, ack => convTransposeC_CP_5782_elements(24)); -- 
    cr_5989_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5989_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(24), ack => RPIPE_Block2_start_2255_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/type_cast_2259_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2255_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2255_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2255_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/type_cast_2259_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2267_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2267_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/type_cast_2259_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2267_sample_start_
      -- 
    ca_5990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2255_inst_ack_1, ack => convTransposeC_CP_5782_elements(25)); -- 
    rr_5998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(25), ack => type_cast_2259_inst_req_0); -- 
    rr_6012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(25), ack => RPIPE_Block2_start_2267_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/type_cast_2259_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/type_cast_2259_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/type_cast_2259_sample_completed_
      -- 
    ra_5999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2259_inst_ack_0, ack => convTransposeC_CP_5782_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/type_cast_2259_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/type_cast_2259_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/type_cast_2259_update_completed_
      -- 
    ca_6004_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2259_inst_ack_1, ack => convTransposeC_CP_5782_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2267_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2267_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2267_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2267_Update/cr
      -- CP-element group 28: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2267_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2267_update_start_
      -- 
    ra_6013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2267_inst_ack_0, ack => convTransposeC_CP_5782_elements(28)); -- 
    cr_6017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(28), ack => RPIPE_Block2_start_2267_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2267_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2270_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2267_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2267_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2270_Sample/rr
      -- CP-element group 29: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2270_Sample/$entry
      -- 
    ca_6018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2267_inst_ack_1, ack => convTransposeC_CP_5782_elements(29)); -- 
    rr_6026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(29), ack => RPIPE_Block2_start_2270_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2270_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2270_update_start_
      -- CP-element group 30: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2270_Update/cr
      -- CP-element group 30: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2270_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2270_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2270_Sample/$exit
      -- 
    ra_6027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2270_inst_ack_0, ack => convTransposeC_CP_5782_elements(30)); -- 
    cr_6031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(30), ack => RPIPE_Block2_start_2270_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2270_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2273_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2273_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2273_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2270_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2270_update_completed_
      -- 
    ca_6032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2270_inst_ack_1, ack => convTransposeC_CP_5782_elements(31)); -- 
    rr_6040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(31), ack => RPIPE_Block2_start_2273_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2273_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2273_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2273_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2273_Update/cr
      -- CP-element group 32: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2273_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2273_update_start_
      -- 
    ra_6041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2273_inst_ack_0, ack => convTransposeC_CP_5782_elements(32)); -- 
    cr_6045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(32), ack => RPIPE_Block2_start_2273_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2273_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2273_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/RPIPE_Block2_start_2273_update_completed_
      -- 
    ca_6046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2273_inst_ack_1, ack => convTransposeC_CP_5782_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34: 	41 
    -- CP-element group 34: 	42 
    -- CP-element group 34:  members (28) 
      -- CP-element group 34: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2306_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2306_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2306_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2310_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2310_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2306_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2310_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2314_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2306_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2314_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2314_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2314_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2310_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/$entry
      -- CP-element group 34: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2310_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2310_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2314_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2314_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2306_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274__exit__
      -- CP-element group 34: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336__entry__
      -- CP-element group 34: 	 branch_block_stmt_2213/assign_stmt_2216_to_assign_stmt_2274/$exit
      -- CP-element group 34: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2318_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2318_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2318_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2318_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2318_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2318_Update/cr
      -- 
    rr_6057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(34), ack => type_cast_2306_inst_req_0); -- 
    cr_6062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(34), ack => type_cast_2306_inst_req_1); -- 
    cr_6090_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6090_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(34), ack => type_cast_2314_inst_req_1); -- 
    cr_6076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(34), ack => type_cast_2310_inst_req_1); -- 
    rr_6071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(34), ack => type_cast_2310_inst_req_0); -- 
    rr_6085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(34), ack => type_cast_2314_inst_req_0); -- 
    rr_6099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(34), ack => type_cast_2318_inst_req_0); -- 
    cr_6104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(34), ack => type_cast_2318_inst_req_1); -- 
    convTransposeC_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(23) & convTransposeC_CP_5782_elements(27) & convTransposeC_CP_5782_elements(33);
      gj_convTransposeC_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2306_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2306_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2306_Sample/ra
      -- 
    ra_6058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2306_inst_ack_0, ack => convTransposeC_CP_5782_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	43 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2306_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2306_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2306_Update/ca
      -- 
    ca_6063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2306_inst_ack_1, ack => convTransposeC_CP_5782_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2310_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2310_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2310_Sample/ra
      -- 
    ra_6072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2310_inst_ack_0, ack => convTransposeC_CP_5782_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	43 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2310_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2310_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2310_Update/ca
      -- 
    ca_6077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2310_inst_ack_1, ack => convTransposeC_CP_5782_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2314_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2314_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2314_Sample/ra
      -- 
    ra_6086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2314_inst_ack_0, ack => convTransposeC_CP_5782_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	43 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2314_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2314_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2314_update_completed_
      -- 
    ca_6091_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2314_inst_ack_1, ack => convTransposeC_CP_5782_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	34 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2318_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2318_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2318_Sample/ra
      -- 
    ra_6100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2318_inst_ack_0, ack => convTransposeC_CP_5782_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	34 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2318_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2318_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/type_cast_2318_Update/ca
      -- 
    ca_6105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2318_inst_ack_1, ack => convTransposeC_CP_5782_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  place  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	36 
    -- CP-element group 43: 	38 
    -- CP-element group 43: 	40 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	79 
    -- CP-element group 43: 	80 
    -- CP-element group 43: 	81 
    -- CP-element group 43: 	82 
    -- CP-element group 43: 	83 
    -- CP-element group 43:  members (18) 
      -- CP-element group 43: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336/$exit
      -- CP-element group 43: 	 branch_block_stmt_2213/assign_stmt_2281_to_assign_stmt_2336__exit__
      -- CP-element group 43: 	 branch_block_stmt_2213/entry_whilex_xbody
      -- CP-element group 43: 	 branch_block_stmt_2213/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 43: 	 branch_block_stmt_2213/entry_whilex_xbody_PhiReq/phi_stmt_2339/$entry
      -- CP-element group 43: 	 branch_block_stmt_2213/entry_whilex_xbody_PhiReq/phi_stmt_2339/phi_stmt_2339_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_2213/entry_whilex_xbody_PhiReq/phi_stmt_2346/$entry
      -- CP-element group 43: 	 branch_block_stmt_2213/entry_whilex_xbody_PhiReq/phi_stmt_2346/phi_stmt_2346_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_2213/entry_whilex_xbody_PhiReq/phi_stmt_2353/$entry
      -- CP-element group 43: 	 branch_block_stmt_2213/entry_whilex_xbody_PhiReq/phi_stmt_2353/phi_stmt_2353_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_2213/entry_whilex_xbody_PhiReq/phi_stmt_2360/$entry
      -- CP-element group 43: 	 branch_block_stmt_2213/entry_whilex_xbody_PhiReq/phi_stmt_2360/phi_stmt_2360_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_2213/entry_whilex_xbody_PhiReq/phi_stmt_2360/phi_stmt_2360_sources/type_cast_2365/$entry
      -- CP-element group 43: 	 branch_block_stmt_2213/entry_whilex_xbody_PhiReq/phi_stmt_2360/phi_stmt_2360_sources/type_cast_2365/SplitProtocol/$entry
      -- CP-element group 43: 	 branch_block_stmt_2213/entry_whilex_xbody_PhiReq/phi_stmt_2360/phi_stmt_2360_sources/type_cast_2365/SplitProtocol/Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_2213/entry_whilex_xbody_PhiReq/phi_stmt_2360/phi_stmt_2360_sources/type_cast_2365/SplitProtocol/Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_2213/entry_whilex_xbody_PhiReq/phi_stmt_2360/phi_stmt_2360_sources/type_cast_2365/SplitProtocol/Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_2213/entry_whilex_xbody_PhiReq/phi_stmt_2360/phi_stmt_2360_sources/type_cast_2365/SplitProtocol/Update/cr
      -- 
    rr_6505_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6505_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(43), ack => type_cast_2365_inst_req_0); -- 
    cr_6510_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6510_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(43), ack => type_cast_2365_inst_req_1); -- 
    convTransposeC_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(36) & convTransposeC_CP_5782_elements(38) & convTransposeC_CP_5782_elements(40) & convTransposeC_CP_5782_elements(42);
      gj_convTransposeC_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	104 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2400_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2400_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2400_Sample/ra
      -- 
    ra_6117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2400_inst_ack_0, ack => convTransposeC_CP_5782_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	104 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	58 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2400_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2400_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2400_Update/ca
      -- 
    ca_6122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2400_inst_ack_1, ack => convTransposeC_CP_5782_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	104 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2404_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2404_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2404_Sample/ra
      -- 
    ra_6131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2404_inst_ack_0, ack => convTransposeC_CP_5782_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	104 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	58 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2404_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2404_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2404_Update/ca
      -- 
    ca_6136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2404_inst_ack_1, ack => convTransposeC_CP_5782_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	104 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2408_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2408_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2408_Sample/ra
      -- 
    ra_6145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2408_inst_ack_0, ack => convTransposeC_CP_5782_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	104 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2408_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2408_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2408_Update/ca
      -- 
    ca_6150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2408_inst_ack_1, ack => convTransposeC_CP_5782_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	104 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2438_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2438_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2438_Sample/ra
      -- 
    ra_6159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2438_inst_ack_0, ack => convTransposeC_CP_5782_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	104 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (16) 
      -- CP-element group 51: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2438_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2438_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2438_Update/ca
      -- CP-element group 51: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2444_index_resized_1
      -- CP-element group 51: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2444_index_scaled_1
      -- CP-element group 51: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2444_index_computed_1
      -- CP-element group 51: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2444_index_resize_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2444_index_resize_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2444_index_resize_1/index_resize_req
      -- CP-element group 51: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2444_index_resize_1/index_resize_ack
      -- CP-element group 51: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2444_index_scale_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2444_index_scale_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2444_index_scale_1/scale_rename_req
      -- CP-element group 51: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2444_index_scale_1/scale_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2444_final_index_sum_regn_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2444_final_index_sum_regn_Sample/req
      -- 
    ca_6164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2438_inst_ack_1, ack => convTransposeC_CP_5782_elements(51)); -- 
    req_6189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(51), ack => array_obj_ref_2444_index_offset_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	68 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2444_final_index_sum_regn_sample_complete
      -- CP-element group 52: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2444_final_index_sum_regn_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2444_final_index_sum_regn_Sample/ack
      -- 
    ack_6190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2444_index_offset_ack_0, ack => convTransposeC_CP_5782_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	104 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (11) 
      -- CP-element group 53: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/addr_of_2445_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2444_root_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2444_offset_calculated
      -- CP-element group 53: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2444_final_index_sum_regn_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2444_final_index_sum_regn_Update/ack
      -- CP-element group 53: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2444_base_plus_offset/$entry
      -- CP-element group 53: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2444_base_plus_offset/$exit
      -- CP-element group 53: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2444_base_plus_offset/sum_rename_req
      -- CP-element group 53: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2444_base_plus_offset/sum_rename_ack
      -- CP-element group 53: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/addr_of_2445_request/$entry
      -- CP-element group 53: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/addr_of_2445_request/req
      -- 
    ack_6195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2444_index_offset_ack_1, ack => convTransposeC_CP_5782_elements(53)); -- 
    req_6204_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6204_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(53), ack => addr_of_2445_final_reg_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/addr_of_2445_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/addr_of_2445_request/$exit
      -- CP-element group 54: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/addr_of_2445_request/ack
      -- 
    ack_6205_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2445_final_reg_ack_0, ack => convTransposeC_CP_5782_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	104 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (24) 
      -- CP-element group 55: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/addr_of_2445_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/addr_of_2445_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/addr_of_2445_complete/ack
      -- CP-element group 55: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2449_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2449_base_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2449_word_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2449_root_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2449_base_address_resized
      -- CP-element group 55: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2449_base_addr_resize/$entry
      -- CP-element group 55: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2449_base_addr_resize/$exit
      -- CP-element group 55: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2449_base_addr_resize/base_resize_req
      -- CP-element group 55: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2449_base_addr_resize/base_resize_ack
      -- CP-element group 55: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2449_base_plus_offset/$entry
      -- CP-element group 55: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2449_base_plus_offset/$exit
      -- CP-element group 55: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2449_base_plus_offset/sum_rename_req
      -- CP-element group 55: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2449_base_plus_offset/sum_rename_ack
      -- CP-element group 55: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2449_word_addrgen/$entry
      -- CP-element group 55: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2449_word_addrgen/$exit
      -- CP-element group 55: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2449_word_addrgen/root_register_req
      -- CP-element group 55: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2449_word_addrgen/root_register_ack
      -- CP-element group 55: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2449_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2449_Sample/word_access_start/$entry
      -- CP-element group 55: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2449_Sample/word_access_start/word_0/$entry
      -- CP-element group 55: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2449_Sample/word_access_start/word_0/rr
      -- 
    ack_6210_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2445_final_reg_ack_1, ack => convTransposeC_CP_5782_elements(55)); -- 
    rr_6243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(55), ack => ptr_deref_2449_load_0_req_0); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (5) 
      -- CP-element group 56: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2449_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2449_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2449_Sample/word_access_start/$exit
      -- CP-element group 56: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2449_Sample/word_access_start/word_0/$exit
      -- CP-element group 56: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2449_Sample/word_access_start/word_0/ra
      -- 
    ra_6244_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2449_load_0_ack_0, ack => convTransposeC_CP_5782_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	104 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (9) 
      -- CP-element group 57: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2449_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2449_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2449_Update/word_access_complete/$exit
      -- CP-element group 57: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2449_Update/word_access_complete/word_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2449_Update/word_access_complete/word_0/ca
      -- CP-element group 57: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2449_Update/ptr_deref_2449_Merge/$entry
      -- CP-element group 57: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2449_Update/ptr_deref_2449_Merge/$exit
      -- CP-element group 57: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2449_Update/ptr_deref_2449_Merge/merge_req
      -- CP-element group 57: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2449_Update/ptr_deref_2449_Merge/merge_ack
      -- 
    ca_6255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2449_load_0_ack_1, ack => convTransposeC_CP_5782_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	45 
    -- CP-element group 58: 	47 
    -- CP-element group 58: 	49 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (13) 
      -- CP-element group 58: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2467_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2467_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2467_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2467_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2467_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2467_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2467_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2467_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2467_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2467_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2467_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2467_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2467_final_index_sum_regn_Sample/req
      -- 
    req_6285_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6285_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(58), ack => array_obj_ref_2467_index_offset_req_0); -- 
    convTransposeC_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(45) & convTransposeC_CP_5782_elements(47) & convTransposeC_CP_5782_elements(49);
      gj_convTransposeC_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	68 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2467_final_index_sum_regn_sample_complete
      -- CP-element group 59: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2467_final_index_sum_regn_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2467_final_index_sum_regn_Sample/ack
      -- 
    ack_6286_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2467_index_offset_ack_0, ack => convTransposeC_CP_5782_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	104 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (11) 
      -- CP-element group 60: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/addr_of_2468_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2467_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2467_offset_calculated
      -- CP-element group 60: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2467_final_index_sum_regn_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2467_final_index_sum_regn_Update/ack
      -- CP-element group 60: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2467_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2467_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2467_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2467_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/addr_of_2468_request/$entry
      -- CP-element group 60: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/addr_of_2468_request/req
      -- 
    ack_6291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2467_index_offset_ack_1, ack => convTransposeC_CP_5782_elements(60)); -- 
    req_6300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(60), ack => addr_of_2468_final_reg_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/addr_of_2468_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/addr_of_2468_request/$exit
      -- CP-element group 61: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/addr_of_2468_request/ack
      -- 
    ack_6301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2468_final_reg_ack_0, ack => convTransposeC_CP_5782_elements(61)); -- 
    -- CP-element group 62:  fork  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	104 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (19) 
      -- CP-element group 62: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/addr_of_2468_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/addr_of_2468_complete/$exit
      -- CP-element group 62: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/addr_of_2468_complete/ack
      -- CP-element group 62: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2471_base_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2471_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2471_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2471_base_address_resized
      -- CP-element group 62: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2471_base_addr_resize/$entry
      -- CP-element group 62: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2471_base_addr_resize/$exit
      -- CP-element group 62: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2471_base_addr_resize/base_resize_req
      -- CP-element group 62: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2471_base_addr_resize/base_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2471_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2471_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2471_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2471_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2471_word_addrgen/$entry
      -- CP-element group 62: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2471_word_addrgen/$exit
      -- CP-element group 62: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2471_word_addrgen/root_register_req
      -- CP-element group 62: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2471_word_addrgen/root_register_ack
      -- 
    ack_6306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2468_final_reg_ack_1, ack => convTransposeC_CP_5782_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2471_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2471_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2471_Sample/ptr_deref_2471_Split/$entry
      -- CP-element group 63: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2471_Sample/ptr_deref_2471_Split/$exit
      -- CP-element group 63: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2471_Sample/ptr_deref_2471_Split/split_req
      -- CP-element group 63: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2471_Sample/ptr_deref_2471_Split/split_ack
      -- CP-element group 63: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2471_Sample/word_access_start/$entry
      -- CP-element group 63: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2471_Sample/word_access_start/word_0/$entry
      -- CP-element group 63: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2471_Sample/word_access_start/word_0/rr
      -- 
    rr_6344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(63), ack => ptr_deref_2471_store_0_req_0); -- 
    convTransposeC_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(57) & convTransposeC_CP_5782_elements(62);
      gj_convTransposeC_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2471_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2471_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2471_Sample/word_access_start/$exit
      -- CP-element group 64: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2471_Sample/word_access_start/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2471_Sample/word_access_start/word_0/ra
      -- 
    ra_6345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2471_store_0_ack_0, ack => convTransposeC_CP_5782_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	104 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	68 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2471_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2471_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2471_Update/word_access_complete/$exit
      -- CP-element group 65: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2471_Update/word_access_complete/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2471_Update/word_access_complete/word_0/ca
      -- 
    ca_6356_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2471_store_0_ack_1, ack => convTransposeC_CP_5782_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	104 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2476_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2476_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2476_Sample/ra
      -- 
    ra_6365_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2476_inst_ack_0, ack => convTransposeC_CP_5782_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	104 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2476_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2476_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2476_Update/ca
      -- 
    ca_6370_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2476_inst_ack_1, ack => convTransposeC_CP_5782_elements(67)); -- 
    -- CP-element group 68:  branch  join  transition  place  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	52 
    -- CP-element group 68: 	59 
    -- CP-element group 68: 	65 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (10) 
      -- CP-element group 68: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488__exit__
      -- CP-element group 68: 	 branch_block_stmt_2213/if_stmt_2489__entry__
      -- CP-element group 68: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/$exit
      -- CP-element group 68: 	 branch_block_stmt_2213/if_stmt_2489_dead_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_2213/if_stmt_2489_eval_test/$entry
      -- CP-element group 68: 	 branch_block_stmt_2213/if_stmt_2489_eval_test/$exit
      -- CP-element group 68: 	 branch_block_stmt_2213/if_stmt_2489_eval_test/branch_req
      -- CP-element group 68: 	 branch_block_stmt_2213/R_cmp_2490_place
      -- CP-element group 68: 	 branch_block_stmt_2213/if_stmt_2489_if_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_2213/if_stmt_2489_else_link/$entry
      -- 
    branch_req_6378_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6378_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(68), ack => if_stmt_2489_branch_req_0); -- 
    convTransposeC_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(52) & convTransposeC_CP_5782_elements(59) & convTransposeC_CP_5782_elements(65) & convTransposeC_CP_5782_elements(67);
      gj_convTransposeC_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	113 
    -- CP-element group 69: 	114 
    -- CP-element group 69: 	116 
    -- CP-element group 69: 	117 
    -- CP-element group 69: 	119 
    -- CP-element group 69: 	120 
    -- CP-element group 69:  members (40) 
      -- CP-element group 69: 	 branch_block_stmt_2213/merge_stmt_2495__exit__
      -- CP-element group 69: 	 branch_block_stmt_2213/assign_stmt_2501__entry__
      -- CP-element group 69: 	 branch_block_stmt_2213/assign_stmt_2501__exit__
      -- CP-element group 69: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133
      -- CP-element group 69: 	 branch_block_stmt_2213/if_stmt_2489_if_link/$exit
      -- CP-element group 69: 	 branch_block_stmt_2213/if_stmt_2489_if_link/if_choice_transition
      -- CP-element group 69: 	 branch_block_stmt_2213/whilex_xbody_ifx_xthen
      -- CP-element group 69: 	 branch_block_stmt_2213/assign_stmt_2501/$entry
      -- CP-element group 69: 	 branch_block_stmt_2213/assign_stmt_2501/$exit
      -- CP-element group 69: 	 branch_block_stmt_2213/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_2213/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 69: 	 branch_block_stmt_2213/merge_stmt_2495_PhiReqMerge
      -- CP-element group 69: 	 branch_block_stmt_2213/merge_stmt_2495_PhiAck/$entry
      -- CP-element group 69: 	 branch_block_stmt_2213/merge_stmt_2495_PhiAck/$exit
      -- CP-element group 69: 	 branch_block_stmt_2213/merge_stmt_2495_PhiAck/dummy
      -- CP-element group 69: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2547/$entry
      -- CP-element group 69: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2547/phi_stmt_2547_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2547/phi_stmt_2547_sources/type_cast_2550/$entry
      -- CP-element group 69: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2547/phi_stmt_2547_sources/type_cast_2550/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2547/phi_stmt_2547_sources/type_cast_2550/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2547/phi_stmt_2547_sources/type_cast_2550/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2547/phi_stmt_2547_sources/type_cast_2550/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2547/phi_stmt_2547_sources/type_cast_2550/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2554/$entry
      -- CP-element group 69: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/type_cast_2559/$entry
      -- CP-element group 69: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/type_cast_2559/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/type_cast_2559/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/type_cast_2559/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/type_cast_2559/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/type_cast_2559/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2560/$entry
      -- CP-element group 69: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2565/$entry
      -- CP-element group 69: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2565/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2565/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2565/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2565/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2565/SplitProtocol/Update/cr
      -- 
    if_choice_transition_6383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2489_branch_ack_1, ack => convTransposeC_CP_5782_elements(69)); -- 
    rr_6715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(69), ack => type_cast_2550_inst_req_0); -- 
    cr_6720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(69), ack => type_cast_2550_inst_req_1); -- 
    rr_6738_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6738_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(69), ack => type_cast_2559_inst_req_0); -- 
    cr_6743_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6743_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(69), ack => type_cast_2559_inst_req_1); -- 
    rr_6761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(69), ack => type_cast_2565_inst_req_0); -- 
    cr_6766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(69), ack => type_cast_2565_inst_req_1); -- 
    -- CP-element group 70:  fork  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70: 	74 
    -- CP-element group 70:  members (21) 
      -- CP-element group 70: 	 branch_block_stmt_2213/merge_stmt_2503__exit__
      -- CP-element group 70: 	 branch_block_stmt_2213/assign_stmt_2509_to_assign_stmt_2539__entry__
      -- CP-element group 70: 	 branch_block_stmt_2213/if_stmt_2489_else_link/$exit
      -- CP-element group 70: 	 branch_block_stmt_2213/if_stmt_2489_else_link/else_choice_transition
      -- CP-element group 70: 	 branch_block_stmt_2213/whilex_xbody_ifx_xelse
      -- CP-element group 70: 	 branch_block_stmt_2213/assign_stmt_2509_to_assign_stmt_2539/$entry
      -- CP-element group 70: 	 branch_block_stmt_2213/assign_stmt_2509_to_assign_stmt_2539/type_cast_2517_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_2213/assign_stmt_2509_to_assign_stmt_2539/type_cast_2517_update_start_
      -- CP-element group 70: 	 branch_block_stmt_2213/assign_stmt_2509_to_assign_stmt_2539/type_cast_2517_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_2213/assign_stmt_2509_to_assign_stmt_2539/type_cast_2517_Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_2213/assign_stmt_2509_to_assign_stmt_2539/type_cast_2517_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_2213/assign_stmt_2509_to_assign_stmt_2539/type_cast_2517_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_2213/assign_stmt_2509_to_assign_stmt_2539/type_cast_2533_update_start_
      -- CP-element group 70: 	 branch_block_stmt_2213/assign_stmt_2509_to_assign_stmt_2539/type_cast_2533_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_2213/assign_stmt_2509_to_assign_stmt_2539/type_cast_2533_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_2213/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_2213/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 70: 	 branch_block_stmt_2213/merge_stmt_2503_PhiReqMerge
      -- CP-element group 70: 	 branch_block_stmt_2213/merge_stmt_2503_PhiAck/$entry
      -- CP-element group 70: 	 branch_block_stmt_2213/merge_stmt_2503_PhiAck/$exit
      -- CP-element group 70: 	 branch_block_stmt_2213/merge_stmt_2503_PhiAck/dummy
      -- 
    else_choice_transition_6387_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2489_branch_ack_0, ack => convTransposeC_CP_5782_elements(70)); -- 
    rr_6403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(70), ack => type_cast_2517_inst_req_0); -- 
    cr_6408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(70), ack => type_cast_2517_inst_req_1); -- 
    cr_6422_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6422_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(70), ack => type_cast_2533_inst_req_1); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_2213/assign_stmt_2509_to_assign_stmt_2539/type_cast_2517_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_2213/assign_stmt_2509_to_assign_stmt_2539/type_cast_2517_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_2213/assign_stmt_2509_to_assign_stmt_2539/type_cast_2517_Sample/ra
      -- 
    ra_6404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2517_inst_ack_0, ack => convTransposeC_CP_5782_elements(71)); -- 
    -- CP-element group 72:  transition  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (6) 
      -- CP-element group 72: 	 branch_block_stmt_2213/assign_stmt_2509_to_assign_stmt_2539/type_cast_2517_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_2213/assign_stmt_2509_to_assign_stmt_2539/type_cast_2517_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_2213/assign_stmt_2509_to_assign_stmt_2539/type_cast_2517_Update/ca
      -- CP-element group 72: 	 branch_block_stmt_2213/assign_stmt_2509_to_assign_stmt_2539/type_cast_2533_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_2213/assign_stmt_2509_to_assign_stmt_2539/type_cast_2533_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_2213/assign_stmt_2509_to_assign_stmt_2539/type_cast_2533_Sample/rr
      -- 
    ca_6409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2517_inst_ack_1, ack => convTransposeC_CP_5782_elements(72)); -- 
    rr_6417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(72), ack => type_cast_2533_inst_req_0); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_2213/assign_stmt_2509_to_assign_stmt_2539/type_cast_2533_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_2213/assign_stmt_2509_to_assign_stmt_2539/type_cast_2533_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_2213/assign_stmt_2509_to_assign_stmt_2539/type_cast_2533_Sample/ra
      -- 
    ra_6418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2533_inst_ack_0, ack => convTransposeC_CP_5782_elements(73)); -- 
    -- CP-element group 74:  branch  transition  place  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	70 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (13) 
      -- CP-element group 74: 	 branch_block_stmt_2213/assign_stmt_2509_to_assign_stmt_2539__exit__
      -- CP-element group 74: 	 branch_block_stmt_2213/if_stmt_2540__entry__
      -- CP-element group 74: 	 branch_block_stmt_2213/assign_stmt_2509_to_assign_stmt_2539/$exit
      -- CP-element group 74: 	 branch_block_stmt_2213/assign_stmt_2509_to_assign_stmt_2539/type_cast_2533_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_2213/assign_stmt_2509_to_assign_stmt_2539/type_cast_2533_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_2213/assign_stmt_2509_to_assign_stmt_2539/type_cast_2533_Update/ca
      -- CP-element group 74: 	 branch_block_stmt_2213/if_stmt_2540_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_2213/if_stmt_2540_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_2213/if_stmt_2540_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_2213/if_stmt_2540_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_2213/R_cmp122_2541_place
      -- CP-element group 74: 	 branch_block_stmt_2213/if_stmt_2540_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_2213/if_stmt_2540_else_link/$entry
      -- 
    ca_6423_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2533_inst_ack_1, ack => convTransposeC_CP_5782_elements(74)); -- 
    branch_req_6431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(74), ack => if_stmt_2540_branch_req_0); -- 
    -- CP-element group 75:  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (15) 
      -- CP-element group 75: 	 branch_block_stmt_2213/merge_stmt_2574__exit__
      -- CP-element group 75: 	 branch_block_stmt_2213/assign_stmt_2579__entry__
      -- CP-element group 75: 	 branch_block_stmt_2213/if_stmt_2540_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_2213/if_stmt_2540_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_2213/ifx_xelse_whilex_xend
      -- CP-element group 75: 	 branch_block_stmt_2213/assign_stmt_2579/$entry
      -- CP-element group 75: 	 branch_block_stmt_2213/assign_stmt_2579/WPIPE_Block2_done_2576_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_2213/assign_stmt_2579/WPIPE_Block2_done_2576_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_2213/assign_stmt_2579/WPIPE_Block2_done_2576_Sample/req
      -- CP-element group 75: 	 branch_block_stmt_2213/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_2213/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_2213/merge_stmt_2574_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_2213/merge_stmt_2574_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_2213/merge_stmt_2574_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_2213/merge_stmt_2574_PhiAck/dummy
      -- 
    if_choice_transition_6436_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2540_branch_ack_1, ack => convTransposeC_CP_5782_elements(75)); -- 
    req_6456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(75), ack => WPIPE_Block2_done_2576_inst_req_0); -- 
    -- CP-element group 76:  fork  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	105 
    -- CP-element group 76: 	106 
    -- CP-element group 76: 	107 
    -- CP-element group 76: 	109 
    -- CP-element group 76: 	110 
    -- CP-element group 76:  members (22) 
      -- CP-element group 76: 	 branch_block_stmt_2213/if_stmt_2540_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_2213/if_stmt_2540_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133
      -- CP-element group 76: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2547/$entry
      -- CP-element group 76: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2547/phi_stmt_2547_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2554/$entry
      -- CP-element group 76: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/type_cast_2557/$entry
      -- CP-element group 76: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/type_cast_2557/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/type_cast_2557/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/type_cast_2557/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/type_cast_2557/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/type_cast_2557/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2560/$entry
      -- CP-element group 76: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2563/$entry
      -- CP-element group 76: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2563/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2563/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2563/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2563/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2563/SplitProtocol/Update/cr
      -- 
    else_choice_transition_6440_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2540_branch_ack_0, ack => convTransposeC_CP_5782_elements(76)); -- 
    rr_6666_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6666_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(76), ack => type_cast_2557_inst_req_0); -- 
    cr_6671_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6671_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(76), ack => type_cast_2557_inst_req_1); -- 
    rr_6689_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6689_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(76), ack => type_cast_2563_inst_req_0); -- 
    cr_6694_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6694_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(76), ack => type_cast_2563_inst_req_1); -- 
    -- CP-element group 77:  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (6) 
      -- CP-element group 77: 	 branch_block_stmt_2213/assign_stmt_2579/WPIPE_Block2_done_2576_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_2213/assign_stmt_2579/WPIPE_Block2_done_2576_update_start_
      -- CP-element group 77: 	 branch_block_stmt_2213/assign_stmt_2579/WPIPE_Block2_done_2576_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_2213/assign_stmt_2579/WPIPE_Block2_done_2576_Sample/ack
      -- CP-element group 77: 	 branch_block_stmt_2213/assign_stmt_2579/WPIPE_Block2_done_2576_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_2213/assign_stmt_2579/WPIPE_Block2_done_2576_Update/req
      -- 
    ack_6457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2576_inst_ack_0, ack => convTransposeC_CP_5782_elements(77)); -- 
    req_6461_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6461_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(77), ack => WPIPE_Block2_done_2576_inst_req_1); -- 
    -- CP-element group 78:  transition  place  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (16) 
      -- CP-element group 78: 	 $exit
      -- CP-element group 78: 	 branch_block_stmt_2213/$exit
      -- CP-element group 78: 	 branch_block_stmt_2213/branch_block_stmt_2213__exit__
      -- CP-element group 78: 	 branch_block_stmt_2213/assign_stmt_2579__exit__
      -- CP-element group 78: 	 branch_block_stmt_2213/return__
      -- CP-element group 78: 	 branch_block_stmt_2213/merge_stmt_2581__exit__
      -- CP-element group 78: 	 branch_block_stmt_2213/assign_stmt_2579/$exit
      -- CP-element group 78: 	 branch_block_stmt_2213/assign_stmt_2579/WPIPE_Block2_done_2576_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_2213/assign_stmt_2579/WPIPE_Block2_done_2576_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_2213/assign_stmt_2579/WPIPE_Block2_done_2576_Update/ack
      -- CP-element group 78: 	 branch_block_stmt_2213/return___PhiReq/$entry
      -- CP-element group 78: 	 branch_block_stmt_2213/return___PhiReq/$exit
      -- CP-element group 78: 	 branch_block_stmt_2213/merge_stmt_2581_PhiReqMerge
      -- CP-element group 78: 	 branch_block_stmt_2213/merge_stmt_2581_PhiAck/$entry
      -- CP-element group 78: 	 branch_block_stmt_2213/merge_stmt_2581_PhiAck/$exit
      -- CP-element group 78: 	 branch_block_stmt_2213/merge_stmt_2581_PhiAck/dummy
      -- 
    ack_6462_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2576_inst_ack_1, ack => convTransposeC_CP_5782_elements(78)); -- 
    -- CP-element group 79:  transition  output  delay-element  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	43 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	85 
    -- CP-element group 79:  members (4) 
      -- CP-element group 79: 	 branch_block_stmt_2213/entry_whilex_xbody_PhiReq/phi_stmt_2339/$exit
      -- CP-element group 79: 	 branch_block_stmt_2213/entry_whilex_xbody_PhiReq/phi_stmt_2339/phi_stmt_2339_sources/$exit
      -- CP-element group 79: 	 branch_block_stmt_2213/entry_whilex_xbody_PhiReq/phi_stmt_2339/phi_stmt_2339_sources/type_cast_2343_konst_delay_trans
      -- CP-element group 79: 	 branch_block_stmt_2213/entry_whilex_xbody_PhiReq/phi_stmt_2339/phi_stmt_2339_req
      -- 
    phi_stmt_2339_req_6473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2339_req_6473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(79), ack => phi_stmt_2339_req_0); -- 
    -- Element group convTransposeC_CP_5782_elements(79) is a control-delay.
    cp_element_79_delay: control_delay_element  generic map(name => " 79_delay", delay_value => 1)  port map(req => convTransposeC_CP_5782_elements(43), ack => convTransposeC_CP_5782_elements(79), clk => clk, reset =>reset);
    -- CP-element group 80:  transition  output  delay-element  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	43 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	85 
    -- CP-element group 80:  members (4) 
      -- CP-element group 80: 	 branch_block_stmt_2213/entry_whilex_xbody_PhiReq/phi_stmt_2346/$exit
      -- CP-element group 80: 	 branch_block_stmt_2213/entry_whilex_xbody_PhiReq/phi_stmt_2346/phi_stmt_2346_sources/$exit
      -- CP-element group 80: 	 branch_block_stmt_2213/entry_whilex_xbody_PhiReq/phi_stmt_2346/phi_stmt_2346_sources/type_cast_2350_konst_delay_trans
      -- CP-element group 80: 	 branch_block_stmt_2213/entry_whilex_xbody_PhiReq/phi_stmt_2346/phi_stmt_2346_req
      -- 
    phi_stmt_2346_req_6481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2346_req_6481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(80), ack => phi_stmt_2346_req_0); -- 
    -- Element group convTransposeC_CP_5782_elements(80) is a control-delay.
    cp_element_80_delay: control_delay_element  generic map(name => " 80_delay", delay_value => 1)  port map(req => convTransposeC_CP_5782_elements(43), ack => convTransposeC_CP_5782_elements(80), clk => clk, reset =>reset);
    -- CP-element group 81:  transition  output  delay-element  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	43 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	85 
    -- CP-element group 81:  members (4) 
      -- CP-element group 81: 	 branch_block_stmt_2213/entry_whilex_xbody_PhiReq/phi_stmt_2353/$exit
      -- CP-element group 81: 	 branch_block_stmt_2213/entry_whilex_xbody_PhiReq/phi_stmt_2353/phi_stmt_2353_sources/$exit
      -- CP-element group 81: 	 branch_block_stmt_2213/entry_whilex_xbody_PhiReq/phi_stmt_2353/phi_stmt_2353_sources/type_cast_2359_konst_delay_trans
      -- CP-element group 81: 	 branch_block_stmt_2213/entry_whilex_xbody_PhiReq/phi_stmt_2353/phi_stmt_2353_req
      -- 
    phi_stmt_2353_req_6489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2353_req_6489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(81), ack => phi_stmt_2353_req_1); -- 
    -- Element group convTransposeC_CP_5782_elements(81) is a control-delay.
    cp_element_81_delay: control_delay_element  generic map(name => " 81_delay", delay_value => 1)  port map(req => convTransposeC_CP_5782_elements(43), ack => convTransposeC_CP_5782_elements(81), clk => clk, reset =>reset);
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	43 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_2213/entry_whilex_xbody_PhiReq/phi_stmt_2360/phi_stmt_2360_sources/type_cast_2365/SplitProtocol/Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_2213/entry_whilex_xbody_PhiReq/phi_stmt_2360/phi_stmt_2360_sources/type_cast_2365/SplitProtocol/Sample/ra
      -- 
    ra_6506_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2365_inst_ack_0, ack => convTransposeC_CP_5782_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	43 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_2213/entry_whilex_xbody_PhiReq/phi_stmt_2360/phi_stmt_2360_sources/type_cast_2365/SplitProtocol/Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_2213/entry_whilex_xbody_PhiReq/phi_stmt_2360/phi_stmt_2360_sources/type_cast_2365/SplitProtocol/Update/ca
      -- 
    ca_6511_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2365_inst_ack_1, ack => convTransposeC_CP_5782_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (5) 
      -- CP-element group 84: 	 branch_block_stmt_2213/entry_whilex_xbody_PhiReq/phi_stmt_2360/$exit
      -- CP-element group 84: 	 branch_block_stmt_2213/entry_whilex_xbody_PhiReq/phi_stmt_2360/phi_stmt_2360_sources/$exit
      -- CP-element group 84: 	 branch_block_stmt_2213/entry_whilex_xbody_PhiReq/phi_stmt_2360/phi_stmt_2360_sources/type_cast_2365/$exit
      -- CP-element group 84: 	 branch_block_stmt_2213/entry_whilex_xbody_PhiReq/phi_stmt_2360/phi_stmt_2360_sources/type_cast_2365/SplitProtocol/$exit
      -- CP-element group 84: 	 branch_block_stmt_2213/entry_whilex_xbody_PhiReq/phi_stmt_2360/phi_stmt_2360_req
      -- 
    phi_stmt_2360_req_6512_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2360_req_6512_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(84), ack => phi_stmt_2360_req_1); -- 
    convTransposeC_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(82) & convTransposeC_CP_5782_elements(83);
      gj_convTransposeC_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  join  transition  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	79 
    -- CP-element group 85: 	80 
    -- CP-element group 85: 	81 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	99 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_2213/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(79) & convTransposeC_CP_5782_elements(80) & convTransposeC_CP_5782_elements(81) & convTransposeC_CP_5782_elements(84);
      gj_convTransposeC_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	1 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2339/phi_stmt_2339_sources/type_cast_2345/SplitProtocol/Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2339/phi_stmt_2339_sources/type_cast_2345/SplitProtocol/Sample/ra
      -- 
    ra_6532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2345_inst_ack_0, ack => convTransposeC_CP_5782_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	1 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2339/phi_stmt_2339_sources/type_cast_2345/SplitProtocol/Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2339/phi_stmt_2339_sources/type_cast_2345/SplitProtocol/Update/ca
      -- 
    ca_6537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2345_inst_ack_1, ack => convTransposeC_CP_5782_elements(87)); -- 
    -- CP-element group 88:  join  transition  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	98 
    -- CP-element group 88:  members (5) 
      -- CP-element group 88: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2339/$exit
      -- CP-element group 88: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2339/phi_stmt_2339_sources/$exit
      -- CP-element group 88: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2339/phi_stmt_2339_sources/type_cast_2345/$exit
      -- CP-element group 88: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2339/phi_stmt_2339_sources/type_cast_2345/SplitProtocol/$exit
      -- CP-element group 88: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2339/phi_stmt_2339_req
      -- 
    phi_stmt_2339_req_6538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2339_req_6538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(88), ack => phi_stmt_2339_req_1); -- 
    convTransposeC_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(86) & convTransposeC_CP_5782_elements(87);
      gj_convTransposeC_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	1 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2346/phi_stmt_2346_sources/type_cast_2352/SplitProtocol/Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2346/phi_stmt_2346_sources/type_cast_2352/SplitProtocol/Sample/ra
      -- 
    ra_6555_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2352_inst_ack_0, ack => convTransposeC_CP_5782_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	1 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2346/phi_stmt_2346_sources/type_cast_2352/SplitProtocol/Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2346/phi_stmt_2346_sources/type_cast_2352/SplitProtocol/Update/ca
      -- 
    ca_6560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2352_inst_ack_1, ack => convTransposeC_CP_5782_elements(90)); -- 
    -- CP-element group 91:  join  transition  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	98 
    -- CP-element group 91:  members (5) 
      -- CP-element group 91: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2346/$exit
      -- CP-element group 91: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2346/phi_stmt_2346_sources/$exit
      -- CP-element group 91: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2346/phi_stmt_2346_sources/type_cast_2352/$exit
      -- CP-element group 91: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2346/phi_stmt_2346_sources/type_cast_2352/SplitProtocol/$exit
      -- CP-element group 91: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2346/phi_stmt_2346_req
      -- 
    phi_stmt_2346_req_6561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2346_req_6561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(91), ack => phi_stmt_2346_req_1); -- 
    convTransposeC_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(89) & convTransposeC_CP_5782_elements(90);
      gj_convTransposeC_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	1 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2353/phi_stmt_2353_sources/type_cast_2356/SplitProtocol/Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2353/phi_stmt_2353_sources/type_cast_2356/SplitProtocol/Sample/ra
      -- 
    ra_6578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2356_inst_ack_0, ack => convTransposeC_CP_5782_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	1 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2353/phi_stmt_2353_sources/type_cast_2356/SplitProtocol/Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2353/phi_stmt_2353_sources/type_cast_2356/SplitProtocol/Update/ca
      -- 
    ca_6583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2356_inst_ack_1, ack => convTransposeC_CP_5782_elements(93)); -- 
    -- CP-element group 94:  join  transition  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	98 
    -- CP-element group 94:  members (5) 
      -- CP-element group 94: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2353/$exit
      -- CP-element group 94: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2353/phi_stmt_2353_sources/$exit
      -- CP-element group 94: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2353/phi_stmt_2353_sources/type_cast_2356/$exit
      -- CP-element group 94: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2353/phi_stmt_2353_sources/type_cast_2356/SplitProtocol/$exit
      -- CP-element group 94: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2353/phi_stmt_2353_req
      -- 
    phi_stmt_2353_req_6584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2353_req_6584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(94), ack => phi_stmt_2353_req_0); -- 
    convTransposeC_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(92) & convTransposeC_CP_5782_elements(93);
      gj_convTransposeC_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	1 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2360/phi_stmt_2360_sources/type_cast_2363/SplitProtocol/Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2360/phi_stmt_2360_sources/type_cast_2363/SplitProtocol/Sample/ra
      -- 
    ra_6601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2363_inst_ack_0, ack => convTransposeC_CP_5782_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	1 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2360/phi_stmt_2360_sources/type_cast_2363/SplitProtocol/Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2360/phi_stmt_2360_sources/type_cast_2363/SplitProtocol/Update/ca
      -- 
    ca_6606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2363_inst_ack_1, ack => convTransposeC_CP_5782_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2360/$exit
      -- CP-element group 97: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2360/phi_stmt_2360_sources/$exit
      -- CP-element group 97: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2360/phi_stmt_2360_sources/type_cast_2363/$exit
      -- CP-element group 97: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2360/phi_stmt_2360_sources/type_cast_2363/SplitProtocol/$exit
      -- CP-element group 97: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2360/phi_stmt_2360_req
      -- 
    phi_stmt_2360_req_6607_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2360_req_6607_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(97), ack => phi_stmt_2360_req_0); -- 
    convTransposeC_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(95) & convTransposeC_CP_5782_elements(96);
      gj_convTransposeC_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	88 
    -- CP-element group 98: 	91 
    -- CP-element group 98: 	94 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_2213/ifx_xend133_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(88) & convTransposeC_CP_5782_elements(91) & convTransposeC_CP_5782_elements(94) & convTransposeC_CP_5782_elements(97);
      gj_convTransposeC_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  merge  fork  transition  place  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	85 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: 	101 
    -- CP-element group 99: 	102 
    -- CP-element group 99: 	103 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_2213/merge_stmt_2338_PhiReqMerge
      -- CP-element group 99: 	 branch_block_stmt_2213/merge_stmt_2338_PhiAck/$entry
      -- 
    convTransposeC_CP_5782_elements(99) <= OrReduce(convTransposeC_CP_5782_elements(85) & convTransposeC_CP_5782_elements(98));
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	104 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_2213/merge_stmt_2338_PhiAck/phi_stmt_2339_ack
      -- 
    phi_stmt_2339_ack_6612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2339_ack_0, ack => convTransposeC_CP_5782_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	104 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_2213/merge_stmt_2338_PhiAck/phi_stmt_2346_ack
      -- 
    phi_stmt_2346_ack_6613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2346_ack_0, ack => convTransposeC_CP_5782_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	99 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_2213/merge_stmt_2338_PhiAck/phi_stmt_2353_ack
      -- 
    phi_stmt_2353_ack_6614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2353_ack_0, ack => convTransposeC_CP_5782_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	99 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_2213/merge_stmt_2338_PhiAck/phi_stmt_2360_ack
      -- 
    phi_stmt_2360_ack_6615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2360_ack_0, ack => convTransposeC_CP_5782_elements(103)); -- 
    -- CP-element group 104:  join  fork  transition  place  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	100 
    -- CP-element group 104: 	101 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	44 
    -- CP-element group 104: 	45 
    -- CP-element group 104: 	46 
    -- CP-element group 104: 	47 
    -- CP-element group 104: 	48 
    -- CP-element group 104: 	49 
    -- CP-element group 104: 	50 
    -- CP-element group 104: 	51 
    -- CP-element group 104: 	53 
    -- CP-element group 104: 	55 
    -- CP-element group 104: 	57 
    -- CP-element group 104: 	60 
    -- CP-element group 104: 	62 
    -- CP-element group 104: 	65 
    -- CP-element group 104: 	66 
    -- CP-element group 104: 	67 
    -- CP-element group 104:  members (56) 
      -- CP-element group 104: 	 branch_block_stmt_2213/merge_stmt_2338__exit__
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488__entry__
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/$entry
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2400_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2400_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2400_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2400_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2400_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2400_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2404_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2404_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2404_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2404_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2404_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2404_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2408_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2408_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2408_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2408_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2408_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2408_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2438_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2438_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2438_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2438_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2438_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2438_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/addr_of_2445_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2444_final_index_sum_regn_update_start
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2444_final_index_sum_regn_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2444_final_index_sum_regn_Update/req
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/addr_of_2445_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/addr_of_2445_complete/req
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2449_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2449_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2449_Update/word_access_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2449_Update/word_access_complete/word_0/$entry
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2449_Update/word_access_complete/word_0/cr
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/addr_of_2468_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2467_final_index_sum_regn_update_start
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2467_final_index_sum_regn_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/array_obj_ref_2467_final_index_sum_regn_Update/req
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/addr_of_2468_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/addr_of_2468_complete/req
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2471_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2471_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2471_Update/word_access_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2471_Update/word_access_complete/word_0/$entry
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/ptr_deref_2471_Update/word_access_complete/word_0/cr
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2476_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2476_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2476_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2476_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2476_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2213/assign_stmt_2372_to_assign_stmt_2488/type_cast_2476_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2213/merge_stmt_2338_PhiAck/$exit
      -- 
    rr_6116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(104), ack => type_cast_2400_inst_req_0); -- 
    cr_6121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(104), ack => type_cast_2400_inst_req_1); -- 
    rr_6130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(104), ack => type_cast_2404_inst_req_0); -- 
    cr_6135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(104), ack => type_cast_2404_inst_req_1); -- 
    rr_6144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(104), ack => type_cast_2408_inst_req_0); -- 
    cr_6149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(104), ack => type_cast_2408_inst_req_1); -- 
    rr_6158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(104), ack => type_cast_2438_inst_req_0); -- 
    cr_6163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(104), ack => type_cast_2438_inst_req_1); -- 
    req_6194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(104), ack => array_obj_ref_2444_index_offset_req_1); -- 
    req_6209_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6209_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(104), ack => addr_of_2445_final_reg_req_1); -- 
    cr_6254_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6254_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(104), ack => ptr_deref_2449_load_0_req_1); -- 
    req_6290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(104), ack => array_obj_ref_2467_index_offset_req_1); -- 
    req_6305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(104), ack => addr_of_2468_final_reg_req_1); -- 
    cr_6355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(104), ack => ptr_deref_2471_store_0_req_1); -- 
    rr_6364_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6364_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(104), ack => type_cast_2476_inst_req_0); -- 
    cr_6369_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6369_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(104), ack => type_cast_2476_inst_req_1); -- 
    convTransposeC_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(100) & convTransposeC_CP_5782_elements(101) & convTransposeC_CP_5782_elements(102) & convTransposeC_CP_5782_elements(103);
      gj_convTransposeC_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  transition  output  delay-element  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	76 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	112 
    -- CP-element group 105:  members (4) 
      -- CP-element group 105: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2547/$exit
      -- CP-element group 105: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2547/phi_stmt_2547_sources/$exit
      -- CP-element group 105: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2547/phi_stmt_2547_sources/type_cast_2553_konst_delay_trans
      -- CP-element group 105: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2547/phi_stmt_2547_req
      -- 
    phi_stmt_2547_req_6650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2547_req_6650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(105), ack => phi_stmt_2547_req_1); -- 
    -- Element group convTransposeC_CP_5782_elements(105) is a control-delay.
    cp_element_105_delay: control_delay_element  generic map(name => " 105_delay", delay_value => 1)  port map(req => convTransposeC_CP_5782_elements(76), ack => convTransposeC_CP_5782_elements(105), clk => clk, reset =>reset);
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	76 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/type_cast_2557/SplitProtocol/Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/type_cast_2557/SplitProtocol/Sample/ra
      -- 
    ra_6667_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2557_inst_ack_0, ack => convTransposeC_CP_5782_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	76 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/type_cast_2557/SplitProtocol/Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/type_cast_2557/SplitProtocol/Update/ca
      -- 
    ca_6672_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2557_inst_ack_1, ack => convTransposeC_CP_5782_elements(107)); -- 
    -- CP-element group 108:  join  transition  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	112 
    -- CP-element group 108:  members (5) 
      -- CP-element group 108: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2554/$exit
      -- CP-element group 108: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/$exit
      -- CP-element group 108: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/type_cast_2557/$exit
      -- CP-element group 108: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/type_cast_2557/SplitProtocol/$exit
      -- CP-element group 108: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2554/phi_stmt_2554_req
      -- 
    phi_stmt_2554_req_6673_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2554_req_6673_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(108), ack => phi_stmt_2554_req_0); -- 
    convTransposeC_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(106) & convTransposeC_CP_5782_elements(107);
      gj_convTransposeC_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	76 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2563/SplitProtocol/Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2563/SplitProtocol/Sample/ra
      -- 
    ra_6690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2563_inst_ack_0, ack => convTransposeC_CP_5782_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	76 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2563/SplitProtocol/Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2563/SplitProtocol/Update/ca
      -- 
    ca_6695_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2563_inst_ack_1, ack => convTransposeC_CP_5782_elements(110)); -- 
    -- CP-element group 111:  join  transition  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (5) 
      -- CP-element group 111: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2560/$exit
      -- CP-element group 111: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/$exit
      -- CP-element group 111: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2563/$exit
      -- CP-element group 111: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2563/SplitProtocol/$exit
      -- CP-element group 111: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_req
      -- 
    phi_stmt_2560_req_6696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2560_req_6696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(111), ack => phi_stmt_2560_req_0); -- 
    convTransposeC_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(109) & convTransposeC_CP_5782_elements(110);
      gj_convTransposeC_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  join  transition  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	105 
    -- CP-element group 112: 	108 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	123 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_2213/ifx_xelse_ifx_xend133_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(105) & convTransposeC_CP_5782_elements(108) & convTransposeC_CP_5782_elements(111);
      gj_convTransposeC_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	69 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2547/phi_stmt_2547_sources/type_cast_2550/SplitProtocol/Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2547/phi_stmt_2547_sources/type_cast_2550/SplitProtocol/Sample/ra
      -- 
    ra_6716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2550_inst_ack_0, ack => convTransposeC_CP_5782_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	69 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (2) 
      -- CP-element group 114: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2547/phi_stmt_2547_sources/type_cast_2550/SplitProtocol/Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2547/phi_stmt_2547_sources/type_cast_2550/SplitProtocol/Update/ca
      -- 
    ca_6721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2550_inst_ack_1, ack => convTransposeC_CP_5782_elements(114)); -- 
    -- CP-element group 115:  join  transition  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	122 
    -- CP-element group 115:  members (5) 
      -- CP-element group 115: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2547/$exit
      -- CP-element group 115: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2547/phi_stmt_2547_sources/$exit
      -- CP-element group 115: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2547/phi_stmt_2547_sources/type_cast_2550/$exit
      -- CP-element group 115: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2547/phi_stmt_2547_sources/type_cast_2550/SplitProtocol/$exit
      -- CP-element group 115: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2547/phi_stmt_2547_req
      -- 
    phi_stmt_2547_req_6722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2547_req_6722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(115), ack => phi_stmt_2547_req_0); -- 
    convTransposeC_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(113) & convTransposeC_CP_5782_elements(114);
      gj_convTransposeC_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	69 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (2) 
      -- CP-element group 116: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/type_cast_2559/SplitProtocol/Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/type_cast_2559/SplitProtocol/Sample/ra
      -- 
    ra_6739_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2559_inst_ack_0, ack => convTransposeC_CP_5782_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	69 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/type_cast_2559/SplitProtocol/Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/type_cast_2559/SplitProtocol/Update/ca
      -- 
    ca_6744_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2559_inst_ack_1, ack => convTransposeC_CP_5782_elements(117)); -- 
    -- CP-element group 118:  join  transition  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	122 
    -- CP-element group 118:  members (5) 
      -- CP-element group 118: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2554/$exit
      -- CP-element group 118: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/$exit
      -- CP-element group 118: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/type_cast_2559/$exit
      -- CP-element group 118: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/type_cast_2559/SplitProtocol/$exit
      -- CP-element group 118: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2554/phi_stmt_2554_req
      -- 
    phi_stmt_2554_req_6745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2554_req_6745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(118), ack => phi_stmt_2554_req_1); -- 
    convTransposeC_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(116) & convTransposeC_CP_5782_elements(117);
      gj_convTransposeC_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	69 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2565/SplitProtocol/Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2565/SplitProtocol/Sample/ra
      -- 
    ra_6762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2565_inst_ack_0, ack => convTransposeC_CP_5782_elements(119)); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	69 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2565/SplitProtocol/Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2565/SplitProtocol/Update/ca
      -- 
    ca_6767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2565_inst_ack_1, ack => convTransposeC_CP_5782_elements(120)); -- 
    -- CP-element group 121:  join  transition  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (5) 
      -- CP-element group 121: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2560/$exit
      -- CP-element group 121: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/$exit
      -- CP-element group 121: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2565/$exit
      -- CP-element group 121: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2565/SplitProtocol/$exit
      -- CP-element group 121: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_req
      -- 
    phi_stmt_2560_req_6768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2560_req_6768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(121), ack => phi_stmt_2560_req_1); -- 
    convTransposeC_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(119) & convTransposeC_CP_5782_elements(120);
      gj_convTransposeC_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  join  transition  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	115 
    -- CP-element group 122: 	118 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_2213/ifx_xthen_ifx_xend133_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(115) & convTransposeC_CP_5782_elements(118) & convTransposeC_CP_5782_elements(121);
      gj_convTransposeC_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  merge  fork  transition  place  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	112 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123: 	125 
    -- CP-element group 123: 	126 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_2213/merge_stmt_2546_PhiReqMerge
      -- CP-element group 123: 	 branch_block_stmt_2213/merge_stmt_2546_PhiAck/$entry
      -- 
    convTransposeC_CP_5782_elements(123) <= OrReduce(convTransposeC_CP_5782_elements(112) & convTransposeC_CP_5782_elements(122));
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	127 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_2213/merge_stmt_2546_PhiAck/phi_stmt_2547_ack
      -- 
    phi_stmt_2547_ack_6773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2547_ack_0, ack => convTransposeC_CP_5782_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_2213/merge_stmt_2546_PhiAck/phi_stmt_2554_ack
      -- 
    phi_stmt_2554_ack_6774_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2554_ack_0, ack => convTransposeC_CP_5782_elements(125)); -- 
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	123 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (1) 
      -- CP-element group 126: 	 branch_block_stmt_2213/merge_stmt_2546_PhiAck/phi_stmt_2560_ack
      -- 
    phi_stmt_2560_ack_6775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2560_ack_0, ack => convTransposeC_CP_5782_elements(126)); -- 
    -- CP-element group 127:  join  transition  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	124 
    -- CP-element group 127: 	125 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	1 
    -- CP-element group 127:  members (1) 
      -- CP-element group 127: 	 branch_block_stmt_2213/merge_stmt_2546_PhiAck/$exit
      -- 
    convTransposeC_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(124) & convTransposeC_CP_5782_elements(125) & convTransposeC_CP_5782_elements(126);
      gj_convTransposeC_cp_element_group_127 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(127), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom86_2466_resized : std_logic_vector(13 downto 0);
    signal R_idxprom86_2466_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2443_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2443_scaled : std_logic_vector(13 downto 0);
    signal add121_2336 : std_logic_vector(31 downto 0);
    signal add45_2287 : std_logic_vector(15 downto 0);
    signal add58_2298 : std_logic_vector(15 downto 0);
    signal add77_2419 : std_logic_vector(63 downto 0);
    signal add79_2429 : std_logic_vector(63 downto 0);
    signal add91_2483 : std_logic_vector(31 downto 0);
    signal add98_2501 : std_logic_vector(15 downto 0);
    signal add_2265 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_2377 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2444_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2444_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2444_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2444_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2444_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2444_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2467_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2467_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2467_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2467_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2467_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2467_root_address : std_logic_vector(13 downto 0);
    signal arrayidx82_2446 : std_logic_vector(31 downto 0);
    signal arrayidx87_2469 : std_logic_vector(31 downto 0);
    signal call11_2234 : std_logic_vector(15 downto 0);
    signal call13_2237 : std_logic_vector(15 downto 0);
    signal call14_2240 : std_logic_vector(15 downto 0);
    signal call15_2243 : std_logic_vector(15 downto 0);
    signal call16_2256 : std_logic_vector(15 downto 0);
    signal call18_2268 : std_logic_vector(15 downto 0);
    signal call1_2219 : std_logic_vector(15 downto 0);
    signal call20_2271 : std_logic_vector(15 downto 0);
    signal call22_2274 : std_logic_vector(15 downto 0);
    signal call3_2222 : std_logic_vector(15 downto 0);
    signal call5_2225 : std_logic_vector(15 downto 0);
    signal call7_2228 : std_logic_vector(15 downto 0);
    signal call9_2231 : std_logic_vector(15 downto 0);
    signal call_2216 : std_logic_vector(15 downto 0);
    signal cmp106_2514 : std_logic_vector(0 downto 0);
    signal cmp122_2539 : std_logic_vector(0 downto 0);
    signal cmp_2488 : std_logic_vector(0 downto 0);
    signal conv112_2534 : std_logic_vector(31 downto 0);
    signal conv115_2319 : std_logic_vector(31 downto 0);
    signal conv17_2260 : std_logic_vector(31 downto 0);
    signal conv65_2401 : std_logic_vector(63 downto 0);
    signal conv68_2307 : std_logic_vector(63 downto 0);
    signal conv70_2405 : std_logic_vector(63 downto 0);
    signal conv73_2311 : std_logic_vector(63 downto 0);
    signal conv75_2409 : std_logic_vector(63 downto 0);
    signal conv90_2477 : std_logic_vector(31 downto 0);
    signal conv94_2315 : std_logic_vector(31 downto 0);
    signal conv_2247 : std_logic_vector(31 downto 0);
    signal idxprom86_2462 : std_logic_vector(63 downto 0);
    signal idxprom_2439 : std_logic_vector(63 downto 0);
    signal inc110_2518 : std_logic_vector(15 downto 0);
    signal inc110x_xinput_dim0x_x2_2523 : std_logic_vector(15 downto 0);
    signal inc_2509 : std_logic_vector(15 downto 0);
    signal indvar_2339 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_2572 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_2560 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_2360 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_2554 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_2353 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2530 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_2547 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2346 : std_logic_vector(15 downto 0);
    signal mul54_2392 : std_logic_vector(15 downto 0);
    signal mul76_2414 : std_logic_vector(63 downto 0);
    signal mul78_2424 : std_logic_vector(63 downto 0);
    signal mul_2382 : std_logic_vector(15 downto 0);
    signal ptr_deref_2449_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2449_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2449_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2449_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2449_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2471_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2471_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2471_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2471_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2471_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2471_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_2253 : std_logic_vector(31 downto 0);
    signal shr116137_2325 : std_logic_vector(31 downto 0);
    signal shr120138_2331 : std_logic_vector(31 downto 0);
    signal shr136_2281 : std_logic_vector(15 downto 0);
    signal shr81_2435 : std_logic_vector(31 downto 0);
    signal shr85_2456 : std_logic_vector(63 downto 0);
    signal sub48_2387 : std_logic_vector(15 downto 0);
    signal sub61_2303 : std_logic_vector(15 downto 0);
    signal sub62_2397 : std_logic_vector(15 downto 0);
    signal sub_2292 : std_logic_vector(15 downto 0);
    signal tmp1_2372 : std_logic_vector(31 downto 0);
    signal tmp83_2450 : std_logic_vector(63 downto 0);
    signal type_cast_2251_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2279_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2285_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2296_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2323_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2329_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2343_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2345_wire : std_logic_vector(31 downto 0);
    signal type_cast_2350_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2352_wire : std_logic_vector(15 downto 0);
    signal type_cast_2356_wire : std_logic_vector(15 downto 0);
    signal type_cast_2359_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2363_wire : std_logic_vector(15 downto 0);
    signal type_cast_2365_wire : std_logic_vector(15 downto 0);
    signal type_cast_2370_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2433_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2454_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2460_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2481_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2499_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2507_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2527_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2550_wire : std_logic_vector(15 downto 0);
    signal type_cast_2553_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2557_wire : std_logic_vector(15 downto 0);
    signal type_cast_2559_wire : std_logic_vector(15 downto 0);
    signal type_cast_2563_wire : std_logic_vector(15 downto 0);
    signal type_cast_2565_wire : std_logic_vector(15 downto 0);
    signal type_cast_2570_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2578_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_2444_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2444_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2444_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2444_resized_base_address <= "00000000000000";
    array_obj_ref_2467_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2467_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2467_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2467_resized_base_address <= "00000000000000";
    ptr_deref_2449_word_offset_0 <= "00000000000000";
    ptr_deref_2471_word_offset_0 <= "00000000000000";
    type_cast_2251_wire_constant <= "00000000000000000000000000010000";
    type_cast_2279_wire_constant <= "0000000000000001";
    type_cast_2285_wire_constant <= "1111111111111111";
    type_cast_2296_wire_constant <= "1111111111111111";
    type_cast_2323_wire_constant <= "00000000000000000000000000000010";
    type_cast_2329_wire_constant <= "00000000000000000000000000000001";
    type_cast_2343_wire_constant <= "00000000000000000000000000000000";
    type_cast_2350_wire_constant <= "0000000000000000";
    type_cast_2359_wire_constant <= "0000000000000000";
    type_cast_2370_wire_constant <= "00000000000000000000000000000100";
    type_cast_2433_wire_constant <= "00000000000000000000000000000010";
    type_cast_2454_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_2460_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_2481_wire_constant <= "00000000000000000000000000000100";
    type_cast_2499_wire_constant <= "0000000000000100";
    type_cast_2507_wire_constant <= "0000000000000001";
    type_cast_2527_wire_constant <= "0000000000000000";
    type_cast_2553_wire_constant <= "0000000000000000";
    type_cast_2570_wire_constant <= "00000000000000000000000000000001";
    type_cast_2578_wire_constant <= "0000000000000001";
    phi_stmt_2339: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2343_wire_constant & type_cast_2345_wire;
      req <= phi_stmt_2339_req_0 & phi_stmt_2339_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2339",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2339_ack_0,
          idata => idata,
          odata => indvar_2339,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2339
    phi_stmt_2346: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2350_wire_constant & type_cast_2352_wire;
      req <= phi_stmt_2346_req_0 & phi_stmt_2346_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2346",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2346_ack_0,
          idata => idata,
          odata => input_dim2x_x1_2346,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2346
    phi_stmt_2353: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2356_wire & type_cast_2359_wire_constant;
      req <= phi_stmt_2353_req_0 & phi_stmt_2353_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2353",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2353_ack_0,
          idata => idata,
          odata => input_dim1x_x1_2353,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2353
    phi_stmt_2360: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2363_wire & type_cast_2365_wire;
      req <= phi_stmt_2360_req_0 & phi_stmt_2360_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2360",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2360_ack_0,
          idata => idata,
          odata => input_dim0x_x2_2360,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2360
    phi_stmt_2547: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2550_wire & type_cast_2553_wire_constant;
      req <= phi_stmt_2547_req_0 & phi_stmt_2547_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2547",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2547_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_2547,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2547
    phi_stmt_2554: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2557_wire & type_cast_2559_wire;
      req <= phi_stmt_2554_req_0 & phi_stmt_2554_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2554",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2554_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_2554,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2554
    phi_stmt_2560: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2563_wire & type_cast_2565_wire;
      req <= phi_stmt_2560_req_0 & phi_stmt_2560_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2560",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2560_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_2560,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2560
    -- flow-through select operator MUX_2529_inst
    input_dim1x_x2_2530 <= type_cast_2527_wire_constant when (cmp106_2514(0) /=  '0') else inc_2509;
    addr_of_2445_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2445_final_reg_req_0;
      addr_of_2445_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2445_final_reg_req_1;
      addr_of_2445_final_reg_ack_1<= rack(0);
      addr_of_2445_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2445_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2444_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx82_2446,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2468_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2468_final_reg_req_0;
      addr_of_2468_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2468_final_reg_req_1;
      addr_of_2468_final_reg_ack_1<= rack(0);
      addr_of_2468_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2468_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2467_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx87_2469,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2246_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2246_inst_req_0;
      type_cast_2246_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2246_inst_req_1;
      type_cast_2246_inst_ack_1<= rack(0);
      type_cast_2246_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2246_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_2243,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_2247,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2259_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2259_inst_req_0;
      type_cast_2259_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2259_inst_req_1;
      type_cast_2259_inst_ack_1<= rack(0);
      type_cast_2259_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2259_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_2256,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_2260,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2306_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2306_inst_req_0;
      type_cast_2306_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2306_inst_req_1;
      type_cast_2306_inst_ack_1<= rack(0);
      type_cast_2306_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2306_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_2274,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv68_2307,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2310_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2310_inst_req_0;
      type_cast_2310_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2310_inst_req_1;
      type_cast_2310_inst_ack_1<= rack(0);
      type_cast_2310_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2310_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_2271,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_2311,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2314_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2314_inst_req_0;
      type_cast_2314_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2314_inst_req_1;
      type_cast_2314_inst_ack_1<= rack(0);
      type_cast_2314_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2314_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_2222,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv94_2315,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2318_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2318_inst_req_0;
      type_cast_2318_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2318_inst_req_1;
      type_cast_2318_inst_ack_1<= rack(0);
      type_cast_2318_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2318_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_2216,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv115_2319,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2345_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2345_inst_req_0;
      type_cast_2345_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2345_inst_req_1;
      type_cast_2345_inst_ack_1<= rack(0);
      type_cast_2345_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2345_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2572,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2345_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2352_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2352_inst_req_0;
      type_cast_2352_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2352_inst_req_1;
      type_cast_2352_inst_ack_1<= rack(0);
      type_cast_2352_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2352_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_2547,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2352_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2356_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2356_inst_req_0;
      type_cast_2356_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2356_inst_req_1;
      type_cast_2356_inst_ack_1<= rack(0);
      type_cast_2356_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2356_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_2554,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2356_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2363_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2363_inst_req_0;
      type_cast_2363_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2363_inst_req_1;
      type_cast_2363_inst_ack_1<= rack(0);
      type_cast_2363_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2363_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_2560,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2363_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2365_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2365_inst_req_0;
      type_cast_2365_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2365_inst_req_1;
      type_cast_2365_inst_ack_1<= rack(0);
      type_cast_2365_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2365_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr136_2281,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2365_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2400_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2400_inst_req_0;
      type_cast_2400_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2400_inst_req_1;
      type_cast_2400_inst_ack_1<= rack(0);
      type_cast_2400_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2400_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2346,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_2401,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2404_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2404_inst_req_0;
      type_cast_2404_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2404_inst_req_1;
      type_cast_2404_inst_ack_1<= rack(0);
      type_cast_2404_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2404_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub62_2397,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_2405,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2408_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2408_inst_req_0;
      type_cast_2408_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2408_inst_req_1;
      type_cast_2408_inst_ack_1<= rack(0);
      type_cast_2408_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2408_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub48_2387,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_2409,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2438_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2438_inst_req_0;
      type_cast_2438_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2438_inst_req_1;
      type_cast_2438_inst_ack_1<= rack(0);
      type_cast_2438_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2438_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr81_2435,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2439,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2476_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2476_inst_req_0;
      type_cast_2476_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2476_inst_req_1;
      type_cast_2476_inst_ack_1<= rack(0);
      type_cast_2476_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2476_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2346,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_2477,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2517_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2517_inst_req_0;
      type_cast_2517_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2517_inst_req_1;
      type_cast_2517_inst_ack_1<= rack(0);
      type_cast_2517_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2517_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp106_2514,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc110_2518,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2533_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2533_inst_req_0;
      type_cast_2533_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2533_inst_req_1;
      type_cast_2533_inst_ack_1<= rack(0);
      type_cast_2533_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2533_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc110x_xinput_dim0x_x2_2523,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv112_2534,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2550_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2550_inst_req_0;
      type_cast_2550_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2550_inst_req_1;
      type_cast_2550_inst_ack_1<= rack(0);
      type_cast_2550_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2550_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add98_2501,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2550_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2557_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2557_inst_req_0;
      type_cast_2557_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2557_inst_req_1;
      type_cast_2557_inst_ack_1<= rack(0);
      type_cast_2557_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2557_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2530,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2557_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2559_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2559_inst_req_0;
      type_cast_2559_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2559_inst_req_1;
      type_cast_2559_inst_ack_1<= rack(0);
      type_cast_2559_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2559_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_2353,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2559_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2563_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2563_inst_req_0;
      type_cast_2563_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2563_inst_req_1;
      type_cast_2563_inst_ack_1<= rack(0);
      type_cast_2563_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2563_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc110x_xinput_dim0x_x2_2523,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2563_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2565_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2565_inst_req_0;
      type_cast_2565_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2565_inst_req_1;
      type_cast_2565_inst_ack_1<= rack(0);
      type_cast_2565_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2565_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_2360,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2565_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_2444_index_1_rename
    process(R_idxprom_2443_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2443_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2443_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2444_index_1_resize
    process(idxprom_2439) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2439;
      ov := iv(13 downto 0);
      R_idxprom_2443_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2444_root_address_inst
    process(array_obj_ref_2444_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2444_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2444_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2467_index_1_rename
    process(R_idxprom86_2466_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom86_2466_resized;
      ov(13 downto 0) := iv;
      R_idxprom86_2466_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2467_index_1_resize
    process(idxprom86_2462) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom86_2462;
      ov := iv(13 downto 0);
      R_idxprom86_2466_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2467_root_address_inst
    process(array_obj_ref_2467_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2467_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2467_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2449_addr_0
    process(ptr_deref_2449_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2449_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2449_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2449_base_resize
    process(arrayidx82_2446) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx82_2446;
      ov := iv(13 downto 0);
      ptr_deref_2449_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2449_gather_scatter
    process(ptr_deref_2449_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2449_data_0;
      ov(63 downto 0) := iv;
      tmp83_2450 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2449_root_address_inst
    process(ptr_deref_2449_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2449_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2449_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2471_addr_0
    process(ptr_deref_2471_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2471_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2471_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2471_base_resize
    process(arrayidx87_2469) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx87_2469;
      ov := iv(13 downto 0);
      ptr_deref_2471_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2471_gather_scatter
    process(tmp83_2450) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp83_2450;
      ov(63 downto 0) := iv;
      ptr_deref_2471_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2471_root_address_inst
    process(ptr_deref_2471_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2471_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2471_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2489_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2488;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2489_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2489_branch_req_0,
          ack0 => if_stmt_2489_branch_ack_0,
          ack1 => if_stmt_2489_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2540_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp122_2539;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2540_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2540_branch_req_0,
          ack0 => if_stmt_2540_branch_ack_0,
          ack1 => if_stmt_2540_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2286_inst
    process(call7_2228) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_2228, type_cast_2285_wire_constant, tmp_var);
      add45_2287 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2297_inst
    process(call9_2231) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_2231, type_cast_2296_wire_constant, tmp_var);
      add58_2298 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2386_inst
    process(sub_2292, mul_2382) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_2292, mul_2382, tmp_var);
      sub48_2387 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2396_inst
    process(sub61_2303, mul54_2392) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub61_2303, mul54_2392, tmp_var);
      sub62_2397 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2500_inst
    process(input_dim2x_x1_2346) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_2346, type_cast_2499_wire_constant, tmp_var);
      add98_2501 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2508_inst
    process(input_dim1x_x1_2353) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_2353, type_cast_2507_wire_constant, tmp_var);
      inc_2509 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2522_inst
    process(inc110_2518, input_dim0x_x2_2360) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc110_2518, input_dim0x_x2_2360, tmp_var);
      inc110x_xinput_dim0x_x2_2523 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2335_inst
    process(shr116137_2325, shr120138_2331) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr116137_2325, shr120138_2331, tmp_var);
      add121_2336 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2376_inst
    process(add_2265, tmp1_2372) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_2265, tmp1_2372, tmp_var);
      add_src_0x_x0_2377 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2482_inst
    process(conv90_2477) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv90_2477, type_cast_2481_wire_constant, tmp_var);
      add91_2483 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2571_inst
    process(indvar_2339) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2339, type_cast_2570_wire_constant, tmp_var);
      indvarx_xnext_2572 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2418_inst
    process(mul76_2414, conv70_2405) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul76_2414, conv70_2405, tmp_var);
      add77_2419 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2428_inst
    process(mul78_2424, conv65_2401) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul78_2424, conv65_2401, tmp_var);
      add79_2429 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2461_inst
    process(shr85_2456) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr85_2456, type_cast_2460_wire_constant, tmp_var);
      idxprom86_2462 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2513_inst
    process(inc_2509, call1_2219) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_2509, call1_2219, tmp_var);
      cmp106_2514 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2538_inst
    process(conv112_2534, add121_2336) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv112_2534, add121_2336, tmp_var);
      cmp122_2539 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2280_inst
    process(call_2216) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_2216, type_cast_2279_wire_constant, tmp_var);
      shr136_2281 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2324_inst
    process(conv115_2319) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv115_2319, type_cast_2323_wire_constant, tmp_var);
      shr116137_2325 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2330_inst
    process(conv115_2319) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv115_2319, type_cast_2329_wire_constant, tmp_var);
      shr120138_2331 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2434_inst
    process(add_src_0x_x0_2377) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_2377, type_cast_2433_wire_constant, tmp_var);
      shr81_2435 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2455_inst
    process(add79_2429) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add79_2429, type_cast_2454_wire_constant, tmp_var);
      shr85_2456 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2381_inst
    process(input_dim0x_x2_2360, call13_2237) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x2_2360, call13_2237, tmp_var);
      mul_2382 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2391_inst
    process(input_dim1x_x1_2353, call13_2237) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_2353, call13_2237, tmp_var);
      mul54_2392 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2371_inst
    process(indvar_2339) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2339, type_cast_2370_wire_constant, tmp_var);
      tmp1_2372 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2413_inst
    process(conv75_2409, conv73_2311) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv75_2409, conv73_2311, tmp_var);
      mul76_2414 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2423_inst
    process(add77_2419, conv68_2307) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add77_2419, conv68_2307, tmp_var);
      mul78_2424 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_2264_inst
    process(shl_2253, conv17_2260) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_2253, conv17_2260, tmp_var);
      add_2265 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2252_inst
    process(conv_2247) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_2247, type_cast_2251_wire_constant, tmp_var);
      shl_2253 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2291_inst
    process(add45_2287, call14_2240) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add45_2287, call14_2240, tmp_var);
      sub_2292 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2302_inst
    process(add58_2298, call14_2240) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add58_2298, call14_2240, tmp_var);
      sub61_2303 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2487_inst
    process(add91_2483, conv94_2315) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add91_2483, conv94_2315, tmp_var);
      cmp_2488 <= tmp_var; --
    end process;
    -- shared split operator group (31) : array_obj_ref_2444_index_offset 
    ApIntAdd_group_31: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2443_scaled;
      array_obj_ref_2444_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2444_index_offset_req_0;
      array_obj_ref_2444_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2444_index_offset_req_1;
      array_obj_ref_2444_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_31_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_31_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_31",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared split operator group (32) : array_obj_ref_2467_index_offset 
    ApIntAdd_group_32: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom86_2466_scaled;
      array_obj_ref_2467_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2467_index_offset_req_0;
      array_obj_ref_2467_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2467_index_offset_req_1;
      array_obj_ref_2467_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_32_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_32_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_32",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- shared load operator group (0) : ptr_deref_2449_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2449_load_0_req_0;
      ptr_deref_2449_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2449_load_0_req_1;
      ptr_deref_2449_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2449_word_address_0;
      ptr_deref_2449_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_2471_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2471_store_0_req_0;
      ptr_deref_2471_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2471_store_0_req_1;
      ptr_deref_2471_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2471_word_address_0;
      data_in <= ptr_deref_2471_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block2_start_2242_inst RPIPE_Block2_start_2255_inst RPIPE_Block2_start_2239_inst RPIPE_Block2_start_2236_inst RPIPE_Block2_start_2233_inst RPIPE_Block2_start_2230_inst RPIPE_Block2_start_2227_inst RPIPE_Block2_start_2224_inst RPIPE_Block2_start_2221_inst RPIPE_Block2_start_2218_inst RPIPE_Block2_start_2273_inst RPIPE_Block2_start_2215_inst RPIPE_Block2_start_2270_inst RPIPE_Block2_start_2267_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block2_start_2242_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block2_start_2255_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block2_start_2239_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block2_start_2236_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block2_start_2233_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block2_start_2230_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block2_start_2227_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block2_start_2224_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block2_start_2221_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block2_start_2218_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block2_start_2273_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block2_start_2215_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block2_start_2270_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block2_start_2267_inst_req_0;
      RPIPE_Block2_start_2242_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block2_start_2255_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block2_start_2239_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block2_start_2236_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block2_start_2233_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block2_start_2230_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block2_start_2227_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block2_start_2224_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block2_start_2221_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block2_start_2218_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block2_start_2273_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block2_start_2215_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block2_start_2270_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block2_start_2267_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block2_start_2242_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block2_start_2255_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block2_start_2239_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block2_start_2236_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block2_start_2233_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block2_start_2230_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block2_start_2227_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block2_start_2224_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block2_start_2221_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block2_start_2218_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block2_start_2273_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block2_start_2215_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block2_start_2270_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block2_start_2267_inst_req_1;
      RPIPE_Block2_start_2242_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block2_start_2255_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block2_start_2239_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block2_start_2236_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block2_start_2233_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block2_start_2230_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block2_start_2227_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block2_start_2224_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block2_start_2221_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block2_start_2218_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block2_start_2273_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block2_start_2215_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block2_start_2270_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block2_start_2267_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call15_2243 <= data_out(223 downto 208);
      call16_2256 <= data_out(207 downto 192);
      call14_2240 <= data_out(191 downto 176);
      call13_2237 <= data_out(175 downto 160);
      call11_2234 <= data_out(159 downto 144);
      call9_2231 <= data_out(143 downto 128);
      call7_2228 <= data_out(127 downto 112);
      call5_2225 <= data_out(111 downto 96);
      call3_2222 <= data_out(95 downto 80);
      call1_2219 <= data_out(79 downto 64);
      call22_2274 <= data_out(63 downto 48);
      call_2216 <= data_out(47 downto 32);
      call20_2271 <= data_out(31 downto 16);
      call18_2268 <= data_out(15 downto 0);
      Block2_start_read_0_gI: SplitGuardInterface generic map(name => "Block2_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_start_read_0: InputPortRevised -- 
        generic map ( name => "Block2_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_start_pipe_read_req(0),
          oack => Block2_start_pipe_read_ack(0),
          odata => Block2_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block2_done_2576_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block2_done_2576_inst_req_0;
      WPIPE_Block2_done_2576_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block2_done_2576_inst_req_1;
      WPIPE_Block2_done_2576_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2578_wire_constant;
      Block2_done_write_0_gI: SplitGuardInterface generic map(name => "Block2_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block2_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_done_pipe_write_req(0),
          oack => Block2_done_pipe_write_ack(0),
          odata => Block2_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeC_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeD is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeD;
architecture convTransposeD_arch of convTransposeD is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeD_CP_6792_start: Boolean;
  signal convTransposeD_CP_6792_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block3_start_2596_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2593_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2614_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2605_inst_req_0 : boolean;
  signal type_cast_2689_inst_req_0 : boolean;
  signal type_cast_2618_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2602_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2596_inst_req_0 : boolean;
  signal type_cast_2766_inst_ack_0 : boolean;
  signal type_cast_2693_inst_req_1 : boolean;
  signal type_cast_2693_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2639_inst_req_1 : boolean;
  signal type_cast_2697_inst_req_0 : boolean;
  signal type_cast_2697_inst_ack_0 : boolean;
  signal type_cast_2618_inst_ack_0 : boolean;
  signal type_cast_2631_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2587_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2602_inst_ack_1 : boolean;
  signal type_cast_2689_inst_req_1 : boolean;
  signal type_cast_2697_inst_req_1 : boolean;
  signal type_cast_2697_inst_ack_1 : boolean;
  signal type_cast_2693_inst_ack_0 : boolean;
  signal type_cast_2762_inst_ack_1 : boolean;
  signal type_cast_2800_inst_req_0 : boolean;
  signal type_cast_2800_inst_ack_0 : boolean;
  signal type_cast_2762_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2602_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2605_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2608_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2587_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2608_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2608_inst_ack_0 : boolean;
  signal type_cast_2631_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2614_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2645_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2639_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2645_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2611_inst_ack_1 : boolean;
  signal type_cast_2618_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2590_inst_ack_1 : boolean;
  signal type_cast_2618_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2596_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2614_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2645_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2602_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2611_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2596_inst_ack_1 : boolean;
  signal type_cast_2631_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2645_inst_ack_0 : boolean;
  signal type_cast_2631_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2593_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2590_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2587_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2614_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2639_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2587_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2642_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2642_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2605_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2642_inst_req_0 : boolean;
  signal type_cast_2689_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2642_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2605_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2590_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2593_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2590_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2639_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2593_inst_ack_1 : boolean;
  signal type_cast_2693_inst_req_0 : boolean;
  signal type_cast_2800_inst_req_1 : boolean;
  signal type_cast_2800_inst_ack_1 : boolean;
  signal type_cast_2762_inst_ack_0 : boolean;
  signal type_cast_2766_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2611_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2611_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2627_inst_ack_1 : boolean;
  signal type_cast_2770_inst_req_0 : boolean;
  signal type_cast_2770_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2627_inst_req_1 : boolean;
  signal array_obj_ref_2806_index_offset_req_0 : boolean;
  signal array_obj_ref_2806_index_offset_ack_0 : boolean;
  signal type_cast_2770_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2599_inst_ack_1 : boolean;
  signal addr_of_2807_final_reg_req_0 : boolean;
  signal addr_of_2807_final_reg_ack_0 : boolean;
  signal addr_of_2807_final_reg_req_1 : boolean;
  signal addr_of_2807_final_reg_ack_1 : boolean;
  signal RPIPE_Block3_start_2599_inst_req_1 : boolean;
  signal array_obj_ref_2806_index_offset_req_1 : boolean;
  signal array_obj_ref_2806_index_offset_ack_1 : boolean;
  signal RPIPE_Block3_start_2599_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2599_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2627_inst_ack_0 : boolean;
  signal type_cast_2770_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2627_inst_req_0 : boolean;
  signal type_cast_2766_inst_req_1 : boolean;
  signal type_cast_2766_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2608_inst_ack_1 : boolean;
  signal type_cast_2762_inst_req_0 : boolean;
  signal type_cast_2689_inst_ack_1 : boolean;
  signal ptr_deref_2811_load_0_req_0 : boolean;
  signal ptr_deref_2811_load_0_ack_0 : boolean;
  signal ptr_deref_2811_load_0_req_1 : boolean;
  signal ptr_deref_2811_load_0_ack_1 : boolean;
  signal array_obj_ref_2829_index_offset_req_0 : boolean;
  signal array_obj_ref_2829_index_offset_ack_0 : boolean;
  signal array_obj_ref_2829_index_offset_req_1 : boolean;
  signal array_obj_ref_2829_index_offset_ack_1 : boolean;
  signal addr_of_2830_final_reg_req_0 : boolean;
  signal addr_of_2830_final_reg_ack_0 : boolean;
  signal addr_of_2830_final_reg_req_1 : boolean;
  signal addr_of_2830_final_reg_ack_1 : boolean;
  signal ptr_deref_2833_store_0_req_0 : boolean;
  signal ptr_deref_2833_store_0_ack_0 : boolean;
  signal ptr_deref_2833_store_0_req_1 : boolean;
  signal ptr_deref_2833_store_0_ack_1 : boolean;
  signal type_cast_2838_inst_req_0 : boolean;
  signal type_cast_2838_inst_ack_0 : boolean;
  signal type_cast_2838_inst_req_1 : boolean;
  signal type_cast_2838_inst_ack_1 : boolean;
  signal if_stmt_2851_branch_req_0 : boolean;
  signal if_stmt_2851_branch_ack_1 : boolean;
  signal if_stmt_2851_branch_ack_0 : boolean;
  signal type_cast_2879_inst_req_0 : boolean;
  signal type_cast_2879_inst_ack_0 : boolean;
  signal type_cast_2879_inst_req_1 : boolean;
  signal type_cast_2879_inst_ack_1 : boolean;
  signal if_stmt_2898_branch_req_0 : boolean;
  signal if_stmt_2898_branch_ack_1 : boolean;
  signal if_stmt_2898_branch_ack_0 : boolean;
  signal WPIPE_Block3_done_2934_inst_req_0 : boolean;
  signal WPIPE_Block3_done_2934_inst_ack_0 : boolean;
  signal WPIPE_Block3_done_2934_inst_req_1 : boolean;
  signal WPIPE_Block3_done_2934_inst_ack_1 : boolean;
  signal phi_stmt_2701_req_0 : boolean;
  signal phi_stmt_2708_req_0 : boolean;
  signal phi_stmt_2715_req_0 : boolean;
  signal type_cast_2725_inst_req_0 : boolean;
  signal type_cast_2725_inst_ack_0 : boolean;
  signal type_cast_2725_inst_req_1 : boolean;
  signal type_cast_2725_inst_ack_1 : boolean;
  signal phi_stmt_2722_req_0 : boolean;
  signal type_cast_2707_inst_req_0 : boolean;
  signal type_cast_2707_inst_ack_0 : boolean;
  signal type_cast_2707_inst_req_1 : boolean;
  signal type_cast_2707_inst_ack_1 : boolean;
  signal phi_stmt_2701_req_1 : boolean;
  signal type_cast_2714_inst_req_0 : boolean;
  signal type_cast_2714_inst_ack_0 : boolean;
  signal type_cast_2714_inst_req_1 : boolean;
  signal type_cast_2714_inst_ack_1 : boolean;
  signal phi_stmt_2708_req_1 : boolean;
  signal type_cast_2721_inst_req_0 : boolean;
  signal type_cast_2721_inst_ack_0 : boolean;
  signal type_cast_2721_inst_req_1 : boolean;
  signal type_cast_2721_inst_ack_1 : boolean;
  signal phi_stmt_2715_req_1 : boolean;
  signal type_cast_2727_inst_req_0 : boolean;
  signal type_cast_2727_inst_ack_0 : boolean;
  signal type_cast_2727_inst_req_1 : boolean;
  signal type_cast_2727_inst_ack_1 : boolean;
  signal phi_stmt_2722_req_1 : boolean;
  signal phi_stmt_2701_ack_0 : boolean;
  signal phi_stmt_2708_ack_0 : boolean;
  signal phi_stmt_2715_ack_0 : boolean;
  signal phi_stmt_2722_ack_0 : boolean;
  signal phi_stmt_2905_req_1 : boolean;
  signal type_cast_2917_inst_req_0 : boolean;
  signal type_cast_2917_inst_ack_0 : boolean;
  signal type_cast_2917_inst_req_1 : boolean;
  signal type_cast_2917_inst_ack_1 : boolean;
  signal phi_stmt_2912_req_1 : boolean;
  signal type_cast_2923_inst_req_0 : boolean;
  signal type_cast_2923_inst_ack_0 : boolean;
  signal type_cast_2923_inst_req_1 : boolean;
  signal type_cast_2923_inst_ack_1 : boolean;
  signal phi_stmt_2918_req_1 : boolean;
  signal type_cast_2908_inst_req_0 : boolean;
  signal type_cast_2908_inst_ack_0 : boolean;
  signal type_cast_2908_inst_req_1 : boolean;
  signal type_cast_2908_inst_ack_1 : boolean;
  signal phi_stmt_2905_req_0 : boolean;
  signal type_cast_2915_inst_req_0 : boolean;
  signal type_cast_2915_inst_ack_0 : boolean;
  signal type_cast_2915_inst_req_1 : boolean;
  signal type_cast_2915_inst_ack_1 : boolean;
  signal phi_stmt_2912_req_0 : boolean;
  signal type_cast_2921_inst_req_0 : boolean;
  signal type_cast_2921_inst_ack_0 : boolean;
  signal type_cast_2921_inst_req_1 : boolean;
  signal type_cast_2921_inst_ack_1 : boolean;
  signal phi_stmt_2918_req_0 : boolean;
  signal phi_stmt_2905_ack_0 : boolean;
  signal phi_stmt_2912_ack_0 : boolean;
  signal phi_stmt_2918_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeD_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeD_CP_6792_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeD_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_6792_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeD_CP_6792_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_6792_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeD_CP_6792: Block -- control-path 
    signal convTransposeD_CP_6792_elements: BooleanArray(123 downto 0);
    -- 
  begin -- 
    convTransposeD_CP_6792_elements(0) <= convTransposeD_CP_6792_start;
    convTransposeD_CP_6792_symbol <= convTransposeD_CP_6792_elements(74);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/type_cast_2631_Update/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2587_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2585/$entry
      -- CP-element group 0: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2587_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/$entry
      -- CP-element group 0: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/type_cast_2618_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/type_cast_2631_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/type_cast_2631_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646__entry__
      -- CP-element group 0: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2587_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/type_cast_2618_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2585/branch_block_stmt_2585__entry__
      -- CP-element group 0: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/type_cast_2618_update_start_
      -- 
    cr_6985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(0), ack => type_cast_2618_inst_req_1); -- 
    cr_7013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(0), ack => type_cast_2631_inst_req_1); -- 
    rr_6840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(0), ack => RPIPE_Block3_start_2587_inst_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	123 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	82 
    -- CP-element group 1: 	83 
    -- CP-element group 1: 	85 
    -- CP-element group 1: 	86 
    -- CP-element group 1: 	88 
    -- CP-element group 1: 	89 
    -- CP-element group 1: 	91 
    -- CP-element group 1: 	92 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_2585/merge_stmt_2904__exit__
      -- CP-element group 1: 	 branch_block_stmt_2585/assign_stmt_2930__exit__
      -- CP-element group 1: 	 branch_block_stmt_2585/assign_stmt_2930__entry__
      -- CP-element group 1: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_2585/assign_stmt_2930/$entry
      -- CP-element group 1: 	 branch_block_stmt_2585/assign_stmt_2930/$exit
      -- CP-element group 1: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2701/$entry
      -- CP-element group 1: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2701/phi_stmt_2701_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2701/phi_stmt_2701_sources/type_cast_2707/$entry
      -- CP-element group 1: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2701/phi_stmt_2701_sources/type_cast_2707/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2701/phi_stmt_2701_sources/type_cast_2707/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2701/phi_stmt_2701_sources/type_cast_2707/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2701/phi_stmt_2701_sources/type_cast_2707/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2701/phi_stmt_2701_sources/type_cast_2707/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2708/$entry
      -- CP-element group 1: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2708/phi_stmt_2708_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2708/phi_stmt_2708_sources/type_cast_2714/$entry
      -- CP-element group 1: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2708/phi_stmt_2708_sources/type_cast_2714/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2708/phi_stmt_2708_sources/type_cast_2714/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2708/phi_stmt_2708_sources/type_cast_2714/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2708/phi_stmt_2708_sources/type_cast_2714/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2708/phi_stmt_2708_sources/type_cast_2714/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2715/$entry
      -- CP-element group 1: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2715/phi_stmt_2715_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2715/phi_stmt_2715_sources/type_cast_2721/$entry
      -- CP-element group 1: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2715/phi_stmt_2715_sources/type_cast_2721/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2715/phi_stmt_2715_sources/type_cast_2721/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2715/phi_stmt_2715_sources/type_cast_2721/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2715/phi_stmt_2715_sources/type_cast_2721/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2715/phi_stmt_2715_sources/type_cast_2721/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2722/$entry
      -- CP-element group 1: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2722/phi_stmt_2722_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2722/phi_stmt_2722_sources/type_cast_2727/$entry
      -- CP-element group 1: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2722/phi_stmt_2722_sources/type_cast_2727/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2722/phi_stmt_2722_sources/type_cast_2727/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2722/phi_stmt_2722_sources/type_cast_2727/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2722/phi_stmt_2722_sources/type_cast_2727/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2722/phi_stmt_2722_sources/type_cast_2727/SplitProtocol/Update/cr
      -- 
    rr_7513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(1), ack => type_cast_2707_inst_req_0); -- 
    cr_7518_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7518_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(1), ack => type_cast_2707_inst_req_1); -- 
    rr_7536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(1), ack => type_cast_2714_inst_req_0); -- 
    cr_7541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(1), ack => type_cast_2714_inst_req_1); -- 
    rr_7559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(1), ack => type_cast_2721_inst_req_0); -- 
    cr_7564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(1), ack => type_cast_2721_inst_req_1); -- 
    rr_7582_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7582_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(1), ack => type_cast_2727_inst_req_0); -- 
    cr_7587_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7587_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(1), ack => type_cast_2727_inst_req_1); -- 
    convTransposeD_CP_6792_elements(1) <= convTransposeD_CP_6792_elements(123);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2587_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2587_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2587_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2587_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2587_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2587_Update/cr
      -- 
    ra_6841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2587_inst_ack_0, ack => convTransposeD_CP_6792_elements(2)); -- 
    cr_6845_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6845_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(2), ack => RPIPE_Block3_start_2587_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2587_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2587_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2587_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2590_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2590_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2590_Sample/rr
      -- 
    ca_6846_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2587_inst_ack_1, ack => convTransposeD_CP_6792_elements(3)); -- 
    rr_6854_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6854_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(3), ack => RPIPE_Block3_start_2590_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2590_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2590_Update/cr
      -- CP-element group 4: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2590_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2590_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2590_update_start_
      -- CP-element group 4: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2590_sample_completed_
      -- 
    ra_6855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2590_inst_ack_0, ack => convTransposeD_CP_6792_elements(4)); -- 
    cr_6859_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6859_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(4), ack => RPIPE_Block3_start_2590_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2593_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2590_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2590_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2593_Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2593_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2590_update_completed_
      -- 
    ca_6860_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2590_inst_ack_1, ack => convTransposeD_CP_6792_elements(5)); -- 
    rr_6868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(5), ack => RPIPE_Block3_start_2593_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2593_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2593_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2593_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2593_update_start_
      -- CP-element group 6: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2593_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2593_Update/cr
      -- 
    ra_6869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2593_inst_ack_0, ack => convTransposeD_CP_6792_elements(6)); -- 
    cr_6873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(6), ack => RPIPE_Block3_start_2593_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2596_Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2593_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2596_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2593_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2593_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2596_sample_start_
      -- 
    ca_6874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2593_inst_ack_1, ack => convTransposeD_CP_6792_elements(7)); -- 
    rr_6882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(7), ack => RPIPE_Block3_start_2596_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2596_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2596_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2596_update_start_
      -- CP-element group 8: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2596_Update/cr
      -- CP-element group 8: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2596_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2596_sample_completed_
      -- 
    ra_6883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2596_inst_ack_0, ack => convTransposeD_CP_6792_elements(8)); -- 
    cr_6887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(8), ack => RPIPE_Block3_start_2596_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2596_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2596_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2596_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2599_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2599_Sample/rr
      -- CP-element group 9: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2599_Sample/$entry
      -- 
    ca_6888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2596_inst_ack_1, ack => convTransposeD_CP_6792_elements(9)); -- 
    rr_6896_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6896_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(9), ack => RPIPE_Block3_start_2599_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2599_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2599_update_start_
      -- CP-element group 10: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2599_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2599_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2599_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2599_Sample/$exit
      -- 
    ra_6897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2599_inst_ack_0, ack => convTransposeD_CP_6792_elements(10)); -- 
    cr_6901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(10), ack => RPIPE_Block3_start_2599_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2602_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2599_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2602_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2602_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2599_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2599_Update/$exit
      -- 
    ca_6902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2599_inst_ack_1, ack => convTransposeD_CP_6792_elements(11)); -- 
    rr_6910_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6910_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(11), ack => RPIPE_Block3_start_2602_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2602_Update/cr
      -- CP-element group 12: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2602_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2602_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2602_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2602_update_start_
      -- CP-element group 12: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2602_sample_completed_
      -- 
    ra_6911_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2602_inst_ack_0, ack => convTransposeD_CP_6792_elements(12)); -- 
    cr_6915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(12), ack => RPIPE_Block3_start_2602_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2605_Sample/rr
      -- CP-element group 13: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2602_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2605_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2602_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2605_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2602_update_completed_
      -- 
    ca_6916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2602_inst_ack_1, ack => convTransposeD_CP_6792_elements(13)); -- 
    rr_6924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(13), ack => RPIPE_Block3_start_2605_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2605_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2605_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2605_update_start_
      -- CP-element group 14: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2605_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2605_Update/cr
      -- CP-element group 14: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2605_Sample/$exit
      -- 
    ra_6925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2605_inst_ack_0, ack => convTransposeD_CP_6792_elements(14)); -- 
    cr_6929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(14), ack => RPIPE_Block3_start_2605_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2605_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2608_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2605_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2605_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2608_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2608_sample_start_
      -- 
    ca_6930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2605_inst_ack_1, ack => convTransposeD_CP_6792_elements(15)); -- 
    rr_6938_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6938_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(15), ack => RPIPE_Block3_start_2608_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2608_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2608_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2608_update_start_
      -- CP-element group 16: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2608_Update/cr
      -- CP-element group 16: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2608_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2608_Update/$entry
      -- 
    ra_6939_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2608_inst_ack_0, ack => convTransposeD_CP_6792_elements(16)); -- 
    cr_6943_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6943_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(16), ack => RPIPE_Block3_start_2608_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2608_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2608_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2611_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2611_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2611_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2608_Update/ca
      -- 
    ca_6944_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2608_inst_ack_1, ack => convTransposeD_CP_6792_elements(17)); -- 
    rr_6952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(17), ack => RPIPE_Block3_start_2611_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2611_Update/cr
      -- CP-element group 18: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2611_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2611_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2611_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2611_update_start_
      -- CP-element group 18: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2611_sample_completed_
      -- 
    ra_6953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2611_inst_ack_0, ack => convTransposeD_CP_6792_elements(18)); -- 
    cr_6957_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6957_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(18), ack => RPIPE_Block3_start_2611_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2611_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2614_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2614_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2611_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2614_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2611_update_completed_
      -- 
    ca_6958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2611_inst_ack_1, ack => convTransposeD_CP_6792_elements(19)); -- 
    rr_6966_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6966_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(19), ack => RPIPE_Block3_start_2614_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2614_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2614_Update/cr
      -- CP-element group 20: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2614_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2614_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2614_update_start_
      -- CP-element group 20: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2614_Sample/$exit
      -- 
    ra_6967_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2614_inst_ack_0, ack => convTransposeD_CP_6792_elements(20)); -- 
    cr_6971_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6971_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(20), ack => RPIPE_Block3_start_2614_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/type_cast_2618_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/type_cast_2618_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2614_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2614_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/type_cast_2618_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2627_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2614_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2627_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2627_Sample/rr
      -- 
    ca_6972_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2614_inst_ack_1, ack => convTransposeD_CP_6792_elements(21)); -- 
    rr_6980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(21), ack => type_cast_2618_inst_req_0); -- 
    rr_6994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(21), ack => RPIPE_Block3_start_2627_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/type_cast_2618_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/type_cast_2618_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/type_cast_2618_sample_completed_
      -- 
    ra_6981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2618_inst_ack_0, ack => convTransposeD_CP_6792_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/type_cast_2618_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/type_cast_2618_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/type_cast_2618_update_completed_
      -- 
    ca_6986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2618_inst_ack_1, ack => convTransposeD_CP_6792_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2627_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2627_update_start_
      -- CP-element group 24: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2627_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2627_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2627_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2627_Sample/$exit
      -- 
    ra_6995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2627_inst_ack_0, ack => convTransposeD_CP_6792_elements(24)); -- 
    cr_6999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(24), ack => RPIPE_Block3_start_2627_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/type_cast_2631_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/type_cast_2631_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2627_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2639_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2639_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2639_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/type_cast_2631_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2627_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2627_Update/$exit
      -- 
    ca_7000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2627_inst_ack_1, ack => convTransposeD_CP_6792_elements(25)); -- 
    rr_7008_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7008_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(25), ack => type_cast_2631_inst_req_0); -- 
    rr_7022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(25), ack => RPIPE_Block3_start_2639_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/type_cast_2631_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/type_cast_2631_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/type_cast_2631_sample_completed_
      -- 
    ra_7009_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2631_inst_ack_0, ack => convTransposeD_CP_6792_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/type_cast_2631_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/type_cast_2631_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/type_cast_2631_Update/ca
      -- 
    ca_7014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2631_inst_ack_1, ack => convTransposeD_CP_6792_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2639_Update/cr
      -- CP-element group 28: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2639_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2639_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2639_update_start_
      -- CP-element group 28: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2639_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2639_Sample/$exit
      -- 
    ra_7023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2639_inst_ack_0, ack => convTransposeD_CP_6792_elements(28)); -- 
    cr_7027_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7027_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(28), ack => RPIPE_Block3_start_2639_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2639_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2642_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2642_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2639_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2642_Sample/rr
      -- CP-element group 29: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2639_update_completed_
      -- 
    ca_7028_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2639_inst_ack_1, ack => convTransposeD_CP_6792_elements(29)); -- 
    rr_7036_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7036_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(29), ack => RPIPE_Block3_start_2642_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2642_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2642_update_start_
      -- CP-element group 30: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2642_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2642_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2642_Update/cr
      -- CP-element group 30: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2642_Sample/ra
      -- 
    ra_7037_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2642_inst_ack_0, ack => convTransposeD_CP_6792_elements(30)); -- 
    cr_7041_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7041_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(30), ack => RPIPE_Block3_start_2642_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2645_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2642_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2642_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2642_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2645_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2645_Sample/$entry
      -- 
    ca_7042_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2642_inst_ack_1, ack => convTransposeD_CP_6792_elements(31)); -- 
    rr_7050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(31), ack => RPIPE_Block3_start_2645_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2645_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2645_Update/cr
      -- CP-element group 32: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2645_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2645_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2645_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2645_update_start_
      -- 
    ra_7051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2645_inst_ack_0, ack => convTransposeD_CP_6792_elements(32)); -- 
    cr_7055_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7055_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(32), ack => RPIPE_Block3_start_2645_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2645_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2645_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/RPIPE_Block3_start_2645_update_completed_
      -- 
    ca_7056_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2645_inst_ack_1, ack => convTransposeD_CP_6792_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34:  members (22) 
      -- CP-element group 34: 	 branch_block_stmt_2585/assign_stmt_2653_to_assign_stmt_2698/type_cast_2689_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2585/assign_stmt_2653_to_assign_stmt_2698/type_cast_2693_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2585/assign_stmt_2653_to_assign_stmt_2698/type_cast_2693_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2585/assign_stmt_2653_to_assign_stmt_2698/type_cast_2697_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2585/assign_stmt_2653_to_assign_stmt_2698/type_cast_2697_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2585/assign_stmt_2653_to_assign_stmt_2698/type_cast_2693_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2585/assign_stmt_2653_to_assign_stmt_2698/type_cast_2693_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2585/assign_stmt_2653_to_assign_stmt_2698/type_cast_2697_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2585/assign_stmt_2653_to_assign_stmt_2698/type_cast_2689_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2585/assign_stmt_2653_to_assign_stmt_2698/type_cast_2689_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646/$exit
      -- CP-element group 34: 	 branch_block_stmt_2585/assign_stmt_2653_to_assign_stmt_2698__entry__
      -- CP-element group 34: 	 branch_block_stmt_2585/assign_stmt_2653_to_assign_stmt_2698/type_cast_2697_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2585/assign_stmt_2653_to_assign_stmt_2698/type_cast_2689_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2585/assign_stmt_2653_to_assign_stmt_2698/type_cast_2697_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2585/assign_stmt_2588_to_assign_stmt_2646__exit__
      -- CP-element group 34: 	 branch_block_stmt_2585/assign_stmt_2653_to_assign_stmt_2698/type_cast_2689_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2585/assign_stmt_2653_to_assign_stmt_2698/type_cast_2697_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2585/assign_stmt_2653_to_assign_stmt_2698/type_cast_2693_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2585/assign_stmt_2653_to_assign_stmt_2698/$entry
      -- CP-element group 34: 	 branch_block_stmt_2585/assign_stmt_2653_to_assign_stmt_2698/type_cast_2693_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2585/assign_stmt_2653_to_assign_stmt_2698/type_cast_2689_update_start_
      -- 
    rr_7067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(34), ack => type_cast_2689_inst_req_0); -- 
    cr_7086_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7086_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(34), ack => type_cast_2693_inst_req_1); -- 
    rr_7095_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7095_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(34), ack => type_cast_2697_inst_req_0); -- 
    cr_7072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(34), ack => type_cast_2689_inst_req_1); -- 
    cr_7100_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7100_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(34), ack => type_cast_2697_inst_req_1); -- 
    rr_7081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(34), ack => type_cast_2693_inst_req_0); -- 
    convTransposeD_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(23) & convTransposeD_CP_6792_elements(27) & convTransposeD_CP_6792_elements(33);
      gj_convTransposeD_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_2585/assign_stmt_2653_to_assign_stmt_2698/type_cast_2689_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_2585/assign_stmt_2653_to_assign_stmt_2698/type_cast_2689_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_2585/assign_stmt_2653_to_assign_stmt_2698/type_cast_2689_Sample/ra
      -- 
    ra_7068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2689_inst_ack_0, ack => convTransposeD_CP_6792_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	41 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_2585/assign_stmt_2653_to_assign_stmt_2698/type_cast_2689_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_2585/assign_stmt_2653_to_assign_stmt_2698/type_cast_2689_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_2585/assign_stmt_2653_to_assign_stmt_2698/type_cast_2689_Update/ca
      -- 
    ca_7073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2689_inst_ack_1, ack => convTransposeD_CP_6792_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_2585/assign_stmt_2653_to_assign_stmt_2698/type_cast_2693_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_2585/assign_stmt_2653_to_assign_stmt_2698/type_cast_2693_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_2585/assign_stmt_2653_to_assign_stmt_2698/type_cast_2693_Sample/$exit
      -- 
    ra_7082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2693_inst_ack_0, ack => convTransposeD_CP_6792_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	41 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_2585/assign_stmt_2653_to_assign_stmt_2698/type_cast_2693_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_2585/assign_stmt_2653_to_assign_stmt_2698/type_cast_2693_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_2585/assign_stmt_2653_to_assign_stmt_2698/type_cast_2693_update_completed_
      -- 
    ca_7087_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2693_inst_ack_1, ack => convTransposeD_CP_6792_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_2585/assign_stmt_2653_to_assign_stmt_2698/type_cast_2697_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_2585/assign_stmt_2653_to_assign_stmt_2698/type_cast_2697_Sample/ra
      -- CP-element group 39: 	 branch_block_stmt_2585/assign_stmt_2653_to_assign_stmt_2698/type_cast_2697_sample_completed_
      -- 
    ra_7096_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2697_inst_ack_0, ack => convTransposeD_CP_6792_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_2585/assign_stmt_2653_to_assign_stmt_2698/type_cast_2697_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_2585/assign_stmt_2653_to_assign_stmt_2698/type_cast_2697_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_2585/assign_stmt_2653_to_assign_stmt_2698/type_cast_2697_Update/$exit
      -- 
    ca_7101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2697_inst_ack_1, ack => convTransposeD_CP_6792_elements(40)); -- 
    -- CP-element group 41:  join  fork  transition  place  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	36 
    -- CP-element group 41: 	38 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	75 
    -- CP-element group 41: 	76 
    -- CP-element group 41: 	77 
    -- CP-element group 41: 	78 
    -- CP-element group 41: 	79 
    -- CP-element group 41:  members (18) 
      -- CP-element group 41: 	 branch_block_stmt_2585/entry_whilex_xbody
      -- CP-element group 41: 	 branch_block_stmt_2585/assign_stmt_2653_to_assign_stmt_2698__exit__
      -- CP-element group 41: 	 branch_block_stmt_2585/assign_stmt_2653_to_assign_stmt_2698/$exit
      -- CP-element group 41: 	 branch_block_stmt_2585/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 41: 	 branch_block_stmt_2585/entry_whilex_xbody_PhiReq/phi_stmt_2701/$entry
      -- CP-element group 41: 	 branch_block_stmt_2585/entry_whilex_xbody_PhiReq/phi_stmt_2701/phi_stmt_2701_sources/$entry
      -- CP-element group 41: 	 branch_block_stmt_2585/entry_whilex_xbody_PhiReq/phi_stmt_2708/$entry
      -- CP-element group 41: 	 branch_block_stmt_2585/entry_whilex_xbody_PhiReq/phi_stmt_2708/phi_stmt_2708_sources/$entry
      -- CP-element group 41: 	 branch_block_stmt_2585/entry_whilex_xbody_PhiReq/phi_stmt_2715/$entry
      -- CP-element group 41: 	 branch_block_stmt_2585/entry_whilex_xbody_PhiReq/phi_stmt_2715/phi_stmt_2715_sources/$entry
      -- CP-element group 41: 	 branch_block_stmt_2585/entry_whilex_xbody_PhiReq/phi_stmt_2722/$entry
      -- CP-element group 41: 	 branch_block_stmt_2585/entry_whilex_xbody_PhiReq/phi_stmt_2722/phi_stmt_2722_sources/$entry
      -- CP-element group 41: 	 branch_block_stmt_2585/entry_whilex_xbody_PhiReq/phi_stmt_2722/phi_stmt_2722_sources/type_cast_2725/$entry
      -- CP-element group 41: 	 branch_block_stmt_2585/entry_whilex_xbody_PhiReq/phi_stmt_2722/phi_stmt_2722_sources/type_cast_2725/SplitProtocol/$entry
      -- CP-element group 41: 	 branch_block_stmt_2585/entry_whilex_xbody_PhiReq/phi_stmt_2722/phi_stmt_2722_sources/type_cast_2725/SplitProtocol/Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_2585/entry_whilex_xbody_PhiReq/phi_stmt_2722/phi_stmt_2722_sources/type_cast_2725/SplitProtocol/Sample/rr
      -- CP-element group 41: 	 branch_block_stmt_2585/entry_whilex_xbody_PhiReq/phi_stmt_2722/phi_stmt_2722_sources/type_cast_2725/SplitProtocol/Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_2585/entry_whilex_xbody_PhiReq/phi_stmt_2722/phi_stmt_2722_sources/type_cast_2725/SplitProtocol/Update/cr
      -- 
    rr_7487_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7487_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(41), ack => type_cast_2725_inst_req_0); -- 
    cr_7492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(41), ack => type_cast_2725_inst_req_1); -- 
    convTransposeD_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(36) & convTransposeD_CP_6792_elements(38) & convTransposeD_CP_6792_elements(40);
      gj_convTransposeD_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	100 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2762_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2762_Sample/ra
      -- CP-element group 42: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2762_Sample/$exit
      -- 
    ra_7113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2762_inst_ack_0, ack => convTransposeD_CP_6792_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	100 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	56 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2762_Update/ca
      -- CP-element group 43: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2762_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2762_update_completed_
      -- 
    ca_7118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2762_inst_ack_1, ack => convTransposeD_CP_6792_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	100 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2766_Sample/ra
      -- CP-element group 44: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2766_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2766_Sample/$exit
      -- 
    ra_7127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2766_inst_ack_0, ack => convTransposeD_CP_6792_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	100 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	56 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2766_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2766_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2766_Update/ca
      -- 
    ca_7132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2766_inst_ack_1, ack => convTransposeD_CP_6792_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	100 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2770_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2770_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2770_Sample/ra
      -- 
    ra_7141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2770_inst_ack_0, ack => convTransposeD_CP_6792_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	100 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	56 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2770_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2770_Update/ca
      -- CP-element group 47: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2770_Update/$exit
      -- 
    ca_7146_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2770_inst_ack_1, ack => convTransposeD_CP_6792_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	100 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2800_Sample/ra
      -- CP-element group 48: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2800_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2800_Sample/$exit
      -- 
    ra_7155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2800_inst_ack_0, ack => convTransposeD_CP_6792_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	100 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (16) 
      -- CP-element group 49: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2800_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2800_Update/ca
      -- CP-element group 49: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2806_final_index_sum_regn_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2806_final_index_sum_regn_Sample/req
      -- CP-element group 49: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2806_index_resized_1
      -- CP-element group 49: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2806_index_scaled_1
      -- CP-element group 49: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2806_index_computed_1
      -- CP-element group 49: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2806_index_scale_1/$entry
      -- CP-element group 49: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2806_index_scale_1/$exit
      -- CP-element group 49: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2806_index_scale_1/scale_rename_req
      -- CP-element group 49: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2806_index_scale_1/scale_rename_ack
      -- CP-element group 49: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2800_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2806_index_resize_1/$entry
      -- CP-element group 49: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2806_index_resize_1/$exit
      -- CP-element group 49: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2806_index_resize_1/index_resize_req
      -- CP-element group 49: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2806_index_resize_1/index_resize_ack
      -- 
    ca_7160_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2800_inst_ack_1, ack => convTransposeD_CP_6792_elements(49)); -- 
    req_7185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(49), ack => array_obj_ref_2806_index_offset_req_0); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	66 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2806_final_index_sum_regn_sample_complete
      -- CP-element group 50: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2806_final_index_sum_regn_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2806_final_index_sum_regn_Sample/ack
      -- 
    ack_7186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2806_index_offset_ack_0, ack => convTransposeD_CP_6792_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	100 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (11) 
      -- CP-element group 51: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/addr_of_2807_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2806_root_address_calculated
      -- CP-element group 51: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2806_offset_calculated
      -- CP-element group 51: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/addr_of_2807_request/$entry
      -- CP-element group 51: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/addr_of_2807_request/req
      -- CP-element group 51: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2806_final_index_sum_regn_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2806_final_index_sum_regn_Update/ack
      -- CP-element group 51: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2806_base_plus_offset/$entry
      -- CP-element group 51: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2806_base_plus_offset/$exit
      -- CP-element group 51: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2806_base_plus_offset/sum_rename_req
      -- CP-element group 51: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2806_base_plus_offset/sum_rename_ack
      -- 
    ack_7191_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2806_index_offset_ack_1, ack => convTransposeD_CP_6792_elements(51)); -- 
    req_7200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(51), ack => addr_of_2807_final_reg_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/addr_of_2807_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/addr_of_2807_request/$exit
      -- CP-element group 52: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/addr_of_2807_request/ack
      -- 
    ack_7201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2807_final_reg_ack_0, ack => convTransposeD_CP_6792_elements(52)); -- 
    -- CP-element group 53:  join  fork  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	100 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (24) 
      -- CP-element group 53: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/addr_of_2807_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/addr_of_2807_complete/$exit
      -- CP-element group 53: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/addr_of_2807_complete/ack
      -- CP-element group 53: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2811_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2811_base_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2811_word_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2811_root_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2811_base_address_resized
      -- CP-element group 53: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2811_base_addr_resize/$entry
      -- CP-element group 53: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2811_base_addr_resize/$exit
      -- CP-element group 53: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2811_base_addr_resize/base_resize_req
      -- CP-element group 53: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2811_base_addr_resize/base_resize_ack
      -- CP-element group 53: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2811_base_plus_offset/$entry
      -- CP-element group 53: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2811_base_plus_offset/$exit
      -- CP-element group 53: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2811_base_plus_offset/sum_rename_req
      -- CP-element group 53: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2811_base_plus_offset/sum_rename_ack
      -- CP-element group 53: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2811_word_addrgen/$entry
      -- CP-element group 53: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2811_word_addrgen/$exit
      -- CP-element group 53: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2811_word_addrgen/root_register_req
      -- CP-element group 53: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2811_word_addrgen/root_register_ack
      -- CP-element group 53: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2811_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2811_Sample/word_access_start/$entry
      -- CP-element group 53: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2811_Sample/word_access_start/word_0/$entry
      -- CP-element group 53: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2811_Sample/word_access_start/word_0/rr
      -- 
    ack_7206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2807_final_reg_ack_1, ack => convTransposeD_CP_6792_elements(53)); -- 
    rr_7239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(53), ack => ptr_deref_2811_load_0_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2811_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2811_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2811_Sample/word_access_start/$exit
      -- CP-element group 54: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2811_Sample/word_access_start/word_0/$exit
      -- CP-element group 54: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2811_Sample/word_access_start/word_0/ra
      -- 
    ra_7240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2811_load_0_ack_0, ack => convTransposeD_CP_6792_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	100 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	61 
    -- CP-element group 55:  members (9) 
      -- CP-element group 55: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2811_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2811_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2811_Update/word_access_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2811_Update/word_access_complete/word_0/$exit
      -- CP-element group 55: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2811_Update/word_access_complete/word_0/ca
      -- CP-element group 55: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2811_Update/ptr_deref_2811_Merge/$entry
      -- CP-element group 55: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2811_Update/ptr_deref_2811_Merge/$exit
      -- CP-element group 55: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2811_Update/ptr_deref_2811_Merge/merge_req
      -- CP-element group 55: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2811_Update/ptr_deref_2811_Merge/merge_ack
      -- 
    ca_7251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2811_load_0_ack_1, ack => convTransposeD_CP_6792_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	43 
    -- CP-element group 56: 	45 
    -- CP-element group 56: 	47 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (13) 
      -- CP-element group 56: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2829_index_scale_1/$entry
      -- CP-element group 56: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2829_index_resized_1
      -- CP-element group 56: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2829_index_scaled_1
      -- CP-element group 56: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2829_index_computed_1
      -- CP-element group 56: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2829_index_resize_1/$entry
      -- CP-element group 56: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2829_index_resize_1/$exit
      -- CP-element group 56: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2829_index_resize_1/index_resize_req
      -- CP-element group 56: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2829_index_resize_1/index_resize_ack
      -- CP-element group 56: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2829_index_scale_1/$exit
      -- CP-element group 56: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2829_index_scale_1/scale_rename_req
      -- CP-element group 56: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2829_index_scale_1/scale_rename_ack
      -- CP-element group 56: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2829_final_index_sum_regn_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2829_final_index_sum_regn_Sample/req
      -- 
    req_7281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(56), ack => array_obj_ref_2829_index_offset_req_0); -- 
    convTransposeD_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(43) & convTransposeD_CP_6792_elements(45) & convTransposeD_CP_6792_elements(47);
      gj_convTransposeD_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	66 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2829_final_index_sum_regn_sample_complete
      -- CP-element group 57: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2829_final_index_sum_regn_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2829_final_index_sum_regn_Sample/ack
      -- 
    ack_7282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2829_index_offset_ack_0, ack => convTransposeD_CP_6792_elements(57)); -- 
    -- CP-element group 58:  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	100 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (11) 
      -- CP-element group 58: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/addr_of_2830_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2829_root_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2829_offset_calculated
      -- CP-element group 58: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2829_final_index_sum_regn_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2829_final_index_sum_regn_Update/ack
      -- CP-element group 58: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2829_base_plus_offset/$entry
      -- CP-element group 58: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2829_base_plus_offset/$exit
      -- CP-element group 58: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2829_base_plus_offset/sum_rename_req
      -- CP-element group 58: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2829_base_plus_offset/sum_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/addr_of_2830_request/$entry
      -- CP-element group 58: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/addr_of_2830_request/req
      -- 
    ack_7287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2829_index_offset_ack_1, ack => convTransposeD_CP_6792_elements(58)); -- 
    req_7296_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7296_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(58), ack => addr_of_2830_final_reg_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/addr_of_2830_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/addr_of_2830_request/$exit
      -- CP-element group 59: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/addr_of_2830_request/ack
      -- 
    ack_7297_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2830_final_reg_ack_0, ack => convTransposeD_CP_6792_elements(59)); -- 
    -- CP-element group 60:  fork  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	100 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (19) 
      -- CP-element group 60: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/addr_of_2830_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/addr_of_2830_complete/$exit
      -- CP-element group 60: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/addr_of_2830_complete/ack
      -- CP-element group 60: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2833_base_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2833_word_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2833_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2833_base_address_resized
      -- CP-element group 60: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2833_base_addr_resize/$entry
      -- CP-element group 60: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2833_base_addr_resize/$exit
      -- CP-element group 60: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2833_base_addr_resize/base_resize_req
      -- CP-element group 60: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2833_base_addr_resize/base_resize_ack
      -- CP-element group 60: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2833_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2833_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2833_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2833_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2833_word_addrgen/$entry
      -- CP-element group 60: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2833_word_addrgen/$exit
      -- CP-element group 60: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2833_word_addrgen/root_register_req
      -- CP-element group 60: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2833_word_addrgen/root_register_ack
      -- 
    ack_7302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2830_final_reg_ack_1, ack => convTransposeD_CP_6792_elements(60)); -- 
    -- CP-element group 61:  join  transition  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	55 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (9) 
      -- CP-element group 61: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2833_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2833_Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2833_Sample/ptr_deref_2833_Split/$entry
      -- CP-element group 61: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2833_Sample/ptr_deref_2833_Split/$exit
      -- CP-element group 61: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2833_Sample/ptr_deref_2833_Split/split_req
      -- CP-element group 61: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2833_Sample/ptr_deref_2833_Split/split_ack
      -- CP-element group 61: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2833_Sample/word_access_start/$entry
      -- CP-element group 61: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2833_Sample/word_access_start/word_0/$entry
      -- CP-element group 61: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2833_Sample/word_access_start/word_0/rr
      -- 
    rr_7340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(61), ack => ptr_deref_2833_store_0_req_0); -- 
    convTransposeD_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(55) & convTransposeD_CP_6792_elements(60);
      gj_convTransposeD_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (5) 
      -- CP-element group 62: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2833_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2833_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2833_Sample/word_access_start/$exit
      -- CP-element group 62: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2833_Sample/word_access_start/word_0/$exit
      -- CP-element group 62: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2833_Sample/word_access_start/word_0/ra
      -- 
    ra_7341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2833_store_0_ack_0, ack => convTransposeD_CP_6792_elements(62)); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	100 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	66 
    -- CP-element group 63:  members (5) 
      -- CP-element group 63: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2833_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2833_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2833_Update/word_access_complete/$exit
      -- CP-element group 63: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2833_Update/word_access_complete/word_0/$exit
      -- CP-element group 63: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2833_Update/word_access_complete/word_0/ca
      -- 
    ca_7352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2833_store_0_ack_1, ack => convTransposeD_CP_6792_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	100 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2838_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2838_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2838_Sample/ra
      -- 
    ra_7361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2838_inst_ack_0, ack => convTransposeD_CP_6792_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	100 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2838_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2838_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2838_Update/ca
      -- 
    ca_7366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2838_inst_ack_1, ack => convTransposeD_CP_6792_elements(65)); -- 
    -- CP-element group 66:  branch  join  transition  place  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	50 
    -- CP-element group 66: 	57 
    -- CP-element group 66: 	63 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (10) 
      -- CP-element group 66: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850__exit__
      -- CP-element group 66: 	 branch_block_stmt_2585/if_stmt_2851__entry__
      -- CP-element group 66: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/$exit
      -- CP-element group 66: 	 branch_block_stmt_2585/if_stmt_2851_dead_link/$entry
      -- CP-element group 66: 	 branch_block_stmt_2585/if_stmt_2851_eval_test/$entry
      -- CP-element group 66: 	 branch_block_stmt_2585/if_stmt_2851_eval_test/$exit
      -- CP-element group 66: 	 branch_block_stmt_2585/if_stmt_2851_eval_test/branch_req
      -- CP-element group 66: 	 branch_block_stmt_2585/R_cmp_2852_place
      -- CP-element group 66: 	 branch_block_stmt_2585/if_stmt_2851_if_link/$entry
      -- CP-element group 66: 	 branch_block_stmt_2585/if_stmt_2851_else_link/$entry
      -- 
    branch_req_7374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(66), ack => if_stmt_2851_branch_req_0); -- 
    convTransposeD_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(50) & convTransposeD_CP_6792_elements(57) & convTransposeD_CP_6792_elements(63) & convTransposeD_CP_6792_elements(65);
      gj_convTransposeD_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	109 
    -- CP-element group 67: 	110 
    -- CP-element group 67: 	112 
    -- CP-element group 67: 	113 
    -- CP-element group 67: 	115 
    -- CP-element group 67: 	116 
    -- CP-element group 67:  members (40) 
      -- CP-element group 67: 	 branch_block_stmt_2585/merge_stmt_2857__exit__
      -- CP-element group 67: 	 branch_block_stmt_2585/assign_stmt_2863__entry__
      -- CP-element group 67: 	 branch_block_stmt_2585/assign_stmt_2863__exit__
      -- CP-element group 67: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132
      -- CP-element group 67: 	 branch_block_stmt_2585/if_stmt_2851_if_link/$exit
      -- CP-element group 67: 	 branch_block_stmt_2585/if_stmt_2851_if_link/if_choice_transition
      -- CP-element group 67: 	 branch_block_stmt_2585/whilex_xbody_ifx_xthen
      -- CP-element group 67: 	 branch_block_stmt_2585/assign_stmt_2863/$entry
      -- CP-element group 67: 	 branch_block_stmt_2585/assign_stmt_2863/$exit
      -- CP-element group 67: 	 branch_block_stmt_2585/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 67: 	 branch_block_stmt_2585/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 67: 	 branch_block_stmt_2585/merge_stmt_2857_PhiReqMerge
      -- CP-element group 67: 	 branch_block_stmt_2585/merge_stmt_2857_PhiAck/$entry
      -- CP-element group 67: 	 branch_block_stmt_2585/merge_stmt_2857_PhiAck/$exit
      -- CP-element group 67: 	 branch_block_stmt_2585/merge_stmt_2857_PhiAck/dummy
      -- CP-element group 67: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/$entry
      -- CP-element group 67: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2905/$entry
      -- CP-element group 67: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2905/phi_stmt_2905_sources/$entry
      -- CP-element group 67: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2905/phi_stmt_2905_sources/type_cast_2908/$entry
      -- CP-element group 67: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2905/phi_stmt_2905_sources/type_cast_2908/SplitProtocol/$entry
      -- CP-element group 67: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2905/phi_stmt_2905_sources/type_cast_2908/SplitProtocol/Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2905/phi_stmt_2905_sources/type_cast_2908/SplitProtocol/Sample/rr
      -- CP-element group 67: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2905/phi_stmt_2905_sources/type_cast_2908/SplitProtocol/Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2905/phi_stmt_2905_sources/type_cast_2908/SplitProtocol/Update/cr
      -- CP-element group 67: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2912/$entry
      -- CP-element group 67: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2912/phi_stmt_2912_sources/$entry
      -- CP-element group 67: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2912/phi_stmt_2912_sources/type_cast_2915/$entry
      -- CP-element group 67: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2912/phi_stmt_2912_sources/type_cast_2915/SplitProtocol/$entry
      -- CP-element group 67: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2912/phi_stmt_2912_sources/type_cast_2915/SplitProtocol/Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2912/phi_stmt_2912_sources/type_cast_2915/SplitProtocol/Sample/rr
      -- CP-element group 67: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2912/phi_stmt_2912_sources/type_cast_2915/SplitProtocol/Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2912/phi_stmt_2912_sources/type_cast_2915/SplitProtocol/Update/cr
      -- CP-element group 67: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2918/$entry
      -- CP-element group 67: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/$entry
      -- CP-element group 67: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2921/$entry
      -- CP-element group 67: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2921/SplitProtocol/$entry
      -- CP-element group 67: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2921/SplitProtocol/Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2921/SplitProtocol/Sample/rr
      -- CP-element group 67: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2921/SplitProtocol/Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2921/SplitProtocol/Update/cr
      -- 
    if_choice_transition_7379_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2851_branch_ack_1, ack => convTransposeD_CP_6792_elements(67)); -- 
    rr_7697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(67), ack => type_cast_2908_inst_req_0); -- 
    cr_7702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(67), ack => type_cast_2908_inst_req_1); -- 
    rr_7720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(67), ack => type_cast_2915_inst_req_0); -- 
    cr_7725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(67), ack => type_cast_2915_inst_req_1); -- 
    rr_7743_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7743_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(67), ack => type_cast_2921_inst_req_0); -- 
    cr_7748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(67), ack => type_cast_2921_inst_req_1); -- 
    -- CP-element group 68:  fork  transition  place  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (18) 
      -- CP-element group 68: 	 branch_block_stmt_2585/merge_stmt_2865__exit__
      -- CP-element group 68: 	 branch_block_stmt_2585/assign_stmt_2871_to_assign_stmt_2897__entry__
      -- CP-element group 68: 	 branch_block_stmt_2585/if_stmt_2851_else_link/$exit
      -- CP-element group 68: 	 branch_block_stmt_2585/if_stmt_2851_else_link/else_choice_transition
      -- CP-element group 68: 	 branch_block_stmt_2585/whilex_xbody_ifx_xelse
      -- CP-element group 68: 	 branch_block_stmt_2585/assign_stmt_2871_to_assign_stmt_2897/$entry
      -- CP-element group 68: 	 branch_block_stmt_2585/assign_stmt_2871_to_assign_stmt_2897/type_cast_2879_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_2585/assign_stmt_2871_to_assign_stmt_2897/type_cast_2879_update_start_
      -- CP-element group 68: 	 branch_block_stmt_2585/assign_stmt_2871_to_assign_stmt_2897/type_cast_2879_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_2585/assign_stmt_2871_to_assign_stmt_2897/type_cast_2879_Sample/rr
      -- CP-element group 68: 	 branch_block_stmt_2585/assign_stmt_2871_to_assign_stmt_2897/type_cast_2879_Update/$entry
      -- CP-element group 68: 	 branch_block_stmt_2585/assign_stmt_2871_to_assign_stmt_2897/type_cast_2879_Update/cr
      -- CP-element group 68: 	 branch_block_stmt_2585/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 68: 	 branch_block_stmt_2585/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 68: 	 branch_block_stmt_2585/merge_stmt_2865_PhiReqMerge
      -- CP-element group 68: 	 branch_block_stmt_2585/merge_stmt_2865_PhiAck/$entry
      -- CP-element group 68: 	 branch_block_stmt_2585/merge_stmt_2865_PhiAck/$exit
      -- CP-element group 68: 	 branch_block_stmt_2585/merge_stmt_2865_PhiAck/dummy
      -- 
    else_choice_transition_7383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2851_branch_ack_0, ack => convTransposeD_CP_6792_elements(68)); -- 
    rr_7399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(68), ack => type_cast_2879_inst_req_0); -- 
    cr_7404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(68), ack => type_cast_2879_inst_req_1); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_2585/assign_stmt_2871_to_assign_stmt_2897/type_cast_2879_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_2585/assign_stmt_2871_to_assign_stmt_2897/type_cast_2879_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_2585/assign_stmt_2871_to_assign_stmt_2897/type_cast_2879_Sample/ra
      -- 
    ra_7400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2879_inst_ack_0, ack => convTransposeD_CP_6792_elements(69)); -- 
    -- CP-element group 70:  branch  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (13) 
      -- CP-element group 70: 	 branch_block_stmt_2585/assign_stmt_2871_to_assign_stmt_2897__exit__
      -- CP-element group 70: 	 branch_block_stmt_2585/if_stmt_2898__entry__
      -- CP-element group 70: 	 branch_block_stmt_2585/assign_stmt_2871_to_assign_stmt_2897/$exit
      -- CP-element group 70: 	 branch_block_stmt_2585/assign_stmt_2871_to_assign_stmt_2897/type_cast_2879_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_2585/assign_stmt_2871_to_assign_stmt_2897/type_cast_2879_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_2585/assign_stmt_2871_to_assign_stmt_2897/type_cast_2879_Update/ca
      -- CP-element group 70: 	 branch_block_stmt_2585/if_stmt_2898_dead_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_2585/if_stmt_2898_eval_test/$entry
      -- CP-element group 70: 	 branch_block_stmt_2585/if_stmt_2898_eval_test/$exit
      -- CP-element group 70: 	 branch_block_stmt_2585/if_stmt_2898_eval_test/branch_req
      -- CP-element group 70: 	 branch_block_stmt_2585/R_cmp121_2899_place
      -- CP-element group 70: 	 branch_block_stmt_2585/if_stmt_2898_if_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_2585/if_stmt_2898_else_link/$entry
      -- 
    ca_7405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2879_inst_ack_1, ack => convTransposeD_CP_6792_elements(70)); -- 
    branch_req_7413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(70), ack => if_stmt_2898_branch_req_0); -- 
    -- CP-element group 71:  transition  place  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (15) 
      -- CP-element group 71: 	 branch_block_stmt_2585/merge_stmt_2932__exit__
      -- CP-element group 71: 	 branch_block_stmt_2585/assign_stmt_2937__entry__
      -- CP-element group 71: 	 branch_block_stmt_2585/if_stmt_2898_if_link/$exit
      -- CP-element group 71: 	 branch_block_stmt_2585/if_stmt_2898_if_link/if_choice_transition
      -- CP-element group 71: 	 branch_block_stmt_2585/ifx_xelse_whilex_xend
      -- CP-element group 71: 	 branch_block_stmt_2585/assign_stmt_2937/$entry
      -- CP-element group 71: 	 branch_block_stmt_2585/assign_stmt_2937/WPIPE_Block3_done_2934_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_2585/assign_stmt_2937/WPIPE_Block3_done_2934_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_2585/assign_stmt_2937/WPIPE_Block3_done_2934_Sample/req
      -- CP-element group 71: 	 branch_block_stmt_2585/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 71: 	 branch_block_stmt_2585/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 71: 	 branch_block_stmt_2585/merge_stmt_2932_PhiReqMerge
      -- CP-element group 71: 	 branch_block_stmt_2585/merge_stmt_2932_PhiAck/$entry
      -- CP-element group 71: 	 branch_block_stmt_2585/merge_stmt_2932_PhiAck/$exit
      -- CP-element group 71: 	 branch_block_stmt_2585/merge_stmt_2932_PhiAck/dummy
      -- 
    if_choice_transition_7418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2898_branch_ack_1, ack => convTransposeD_CP_6792_elements(71)); -- 
    req_7438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(71), ack => WPIPE_Block3_done_2934_inst_req_0); -- 
    -- CP-element group 72:  fork  transition  place  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	101 
    -- CP-element group 72: 	102 
    -- CP-element group 72: 	103 
    -- CP-element group 72: 	105 
    -- CP-element group 72: 	106 
    -- CP-element group 72:  members (22) 
      -- CP-element group 72: 	 branch_block_stmt_2585/if_stmt_2898_else_link/$exit
      -- CP-element group 72: 	 branch_block_stmt_2585/if_stmt_2898_else_link/else_choice_transition
      -- CP-element group 72: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132
      -- CP-element group 72: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/$entry
      -- CP-element group 72: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2905/$entry
      -- CP-element group 72: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2905/phi_stmt_2905_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2912/$entry
      -- CP-element group 72: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2912/phi_stmt_2912_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2912/phi_stmt_2912_sources/type_cast_2917/$entry
      -- CP-element group 72: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2912/phi_stmt_2912_sources/type_cast_2917/SplitProtocol/$entry
      -- CP-element group 72: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2912/phi_stmt_2912_sources/type_cast_2917/SplitProtocol/Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2912/phi_stmt_2912_sources/type_cast_2917/SplitProtocol/Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2912/phi_stmt_2912_sources/type_cast_2917/SplitProtocol/Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2912/phi_stmt_2912_sources/type_cast_2917/SplitProtocol/Update/cr
      -- CP-element group 72: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2918/$entry
      -- CP-element group 72: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2923/$entry
      -- CP-element group 72: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2923/SplitProtocol/$entry
      -- CP-element group 72: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2923/SplitProtocol/Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2923/SplitProtocol/Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2923/SplitProtocol/Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2923/SplitProtocol/Update/cr
      -- 
    else_choice_transition_7422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2898_branch_ack_0, ack => convTransposeD_CP_6792_elements(72)); -- 
    rr_7648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(72), ack => type_cast_2917_inst_req_0); -- 
    cr_7653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(72), ack => type_cast_2917_inst_req_1); -- 
    rr_7671_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7671_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(72), ack => type_cast_2923_inst_req_0); -- 
    cr_7676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(72), ack => type_cast_2923_inst_req_1); -- 
    -- CP-element group 73:  transition  input  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (6) 
      -- CP-element group 73: 	 branch_block_stmt_2585/assign_stmt_2937/WPIPE_Block3_done_2934_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_2585/assign_stmt_2937/WPIPE_Block3_done_2934_update_start_
      -- CP-element group 73: 	 branch_block_stmt_2585/assign_stmt_2937/WPIPE_Block3_done_2934_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_2585/assign_stmt_2937/WPIPE_Block3_done_2934_Sample/ack
      -- CP-element group 73: 	 branch_block_stmt_2585/assign_stmt_2937/WPIPE_Block3_done_2934_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_2585/assign_stmt_2937/WPIPE_Block3_done_2934_Update/req
      -- 
    ack_7439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_2934_inst_ack_0, ack => convTransposeD_CP_6792_elements(73)); -- 
    req_7443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(73), ack => WPIPE_Block3_done_2934_inst_req_1); -- 
    -- CP-element group 74:  transition  place  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (16) 
      -- CP-element group 74: 	 $exit
      -- CP-element group 74: 	 branch_block_stmt_2585/merge_stmt_2939__exit__
      -- CP-element group 74: 	 branch_block_stmt_2585/$exit
      -- CP-element group 74: 	 branch_block_stmt_2585/branch_block_stmt_2585__exit__
      -- CP-element group 74: 	 branch_block_stmt_2585/assign_stmt_2937__exit__
      -- CP-element group 74: 	 branch_block_stmt_2585/return__
      -- CP-element group 74: 	 branch_block_stmt_2585/assign_stmt_2937/$exit
      -- CP-element group 74: 	 branch_block_stmt_2585/assign_stmt_2937/WPIPE_Block3_done_2934_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_2585/assign_stmt_2937/WPIPE_Block3_done_2934_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_2585/assign_stmt_2937/WPIPE_Block3_done_2934_Update/ack
      -- CP-element group 74: 	 branch_block_stmt_2585/return___PhiReq/$entry
      -- CP-element group 74: 	 branch_block_stmt_2585/return___PhiReq/$exit
      -- CP-element group 74: 	 branch_block_stmt_2585/merge_stmt_2939_PhiReqMerge
      -- CP-element group 74: 	 branch_block_stmt_2585/merge_stmt_2939_PhiAck/$entry
      -- CP-element group 74: 	 branch_block_stmt_2585/merge_stmt_2939_PhiAck/$exit
      -- CP-element group 74: 	 branch_block_stmt_2585/merge_stmt_2939_PhiAck/dummy
      -- 
    ack_7444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_2934_inst_ack_1, ack => convTransposeD_CP_6792_elements(74)); -- 
    -- CP-element group 75:  transition  output  delay-element  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	41 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	81 
    -- CP-element group 75:  members (4) 
      -- CP-element group 75: 	 branch_block_stmt_2585/entry_whilex_xbody_PhiReq/phi_stmt_2701/$exit
      -- CP-element group 75: 	 branch_block_stmt_2585/entry_whilex_xbody_PhiReq/phi_stmt_2701/phi_stmt_2701_sources/$exit
      -- CP-element group 75: 	 branch_block_stmt_2585/entry_whilex_xbody_PhiReq/phi_stmt_2701/phi_stmt_2701_sources/type_cast_2705_konst_delay_trans
      -- CP-element group 75: 	 branch_block_stmt_2585/entry_whilex_xbody_PhiReq/phi_stmt_2701/phi_stmt_2701_req
      -- 
    phi_stmt_2701_req_7455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2701_req_7455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(75), ack => phi_stmt_2701_req_0); -- 
    -- Element group convTransposeD_CP_6792_elements(75) is a control-delay.
    cp_element_75_delay: control_delay_element  generic map(name => " 75_delay", delay_value => 1)  port map(req => convTransposeD_CP_6792_elements(41), ack => convTransposeD_CP_6792_elements(75), clk => clk, reset =>reset);
    -- CP-element group 76:  transition  output  delay-element  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	41 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	81 
    -- CP-element group 76:  members (4) 
      -- CP-element group 76: 	 branch_block_stmt_2585/entry_whilex_xbody_PhiReq/phi_stmt_2708/$exit
      -- CP-element group 76: 	 branch_block_stmt_2585/entry_whilex_xbody_PhiReq/phi_stmt_2708/phi_stmt_2708_sources/$exit
      -- CP-element group 76: 	 branch_block_stmt_2585/entry_whilex_xbody_PhiReq/phi_stmt_2708/phi_stmt_2708_sources/type_cast_2712_konst_delay_trans
      -- CP-element group 76: 	 branch_block_stmt_2585/entry_whilex_xbody_PhiReq/phi_stmt_2708/phi_stmt_2708_req
      -- 
    phi_stmt_2708_req_7463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2708_req_7463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(76), ack => phi_stmt_2708_req_0); -- 
    -- Element group convTransposeD_CP_6792_elements(76) is a control-delay.
    cp_element_76_delay: control_delay_element  generic map(name => " 76_delay", delay_value => 1)  port map(req => convTransposeD_CP_6792_elements(41), ack => convTransposeD_CP_6792_elements(76), clk => clk, reset =>reset);
    -- CP-element group 77:  transition  output  delay-element  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	41 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	81 
    -- CP-element group 77:  members (4) 
      -- CP-element group 77: 	 branch_block_stmt_2585/entry_whilex_xbody_PhiReq/phi_stmt_2715/$exit
      -- CP-element group 77: 	 branch_block_stmt_2585/entry_whilex_xbody_PhiReq/phi_stmt_2715/phi_stmt_2715_sources/$exit
      -- CP-element group 77: 	 branch_block_stmt_2585/entry_whilex_xbody_PhiReq/phi_stmt_2715/phi_stmt_2715_sources/type_cast_2719_konst_delay_trans
      -- CP-element group 77: 	 branch_block_stmt_2585/entry_whilex_xbody_PhiReq/phi_stmt_2715/phi_stmt_2715_req
      -- 
    phi_stmt_2715_req_7471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2715_req_7471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(77), ack => phi_stmt_2715_req_0); -- 
    -- Element group convTransposeD_CP_6792_elements(77) is a control-delay.
    cp_element_77_delay: control_delay_element  generic map(name => " 77_delay", delay_value => 1)  port map(req => convTransposeD_CP_6792_elements(41), ack => convTransposeD_CP_6792_elements(77), clk => clk, reset =>reset);
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	41 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (2) 
      -- CP-element group 78: 	 branch_block_stmt_2585/entry_whilex_xbody_PhiReq/phi_stmt_2722/phi_stmt_2722_sources/type_cast_2725/SplitProtocol/Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_2585/entry_whilex_xbody_PhiReq/phi_stmt_2722/phi_stmt_2722_sources/type_cast_2725/SplitProtocol/Sample/ra
      -- 
    ra_7488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2725_inst_ack_0, ack => convTransposeD_CP_6792_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	41 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_2585/entry_whilex_xbody_PhiReq/phi_stmt_2722/phi_stmt_2722_sources/type_cast_2725/SplitProtocol/Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_2585/entry_whilex_xbody_PhiReq/phi_stmt_2722/phi_stmt_2722_sources/type_cast_2725/SplitProtocol/Update/ca
      -- 
    ca_7493_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2725_inst_ack_1, ack => convTransposeD_CP_6792_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (5) 
      -- CP-element group 80: 	 branch_block_stmt_2585/entry_whilex_xbody_PhiReq/phi_stmt_2722/$exit
      -- CP-element group 80: 	 branch_block_stmt_2585/entry_whilex_xbody_PhiReq/phi_stmt_2722/phi_stmt_2722_sources/$exit
      -- CP-element group 80: 	 branch_block_stmt_2585/entry_whilex_xbody_PhiReq/phi_stmt_2722/phi_stmt_2722_sources/type_cast_2725/$exit
      -- CP-element group 80: 	 branch_block_stmt_2585/entry_whilex_xbody_PhiReq/phi_stmt_2722/phi_stmt_2722_sources/type_cast_2725/SplitProtocol/$exit
      -- CP-element group 80: 	 branch_block_stmt_2585/entry_whilex_xbody_PhiReq/phi_stmt_2722/phi_stmt_2722_req
      -- 
    phi_stmt_2722_req_7494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2722_req_7494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(80), ack => phi_stmt_2722_req_0); -- 
    convTransposeD_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(78) & convTransposeD_CP_6792_elements(79);
      gj_convTransposeD_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  join  transition  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	75 
    -- CP-element group 81: 	76 
    -- CP-element group 81: 	77 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	95 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_2585/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(75) & convTransposeD_CP_6792_elements(76) & convTransposeD_CP_6792_elements(77) & convTransposeD_CP_6792_elements(80);
      gj_convTransposeD_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	1 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2701/phi_stmt_2701_sources/type_cast_2707/SplitProtocol/Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2701/phi_stmt_2701_sources/type_cast_2707/SplitProtocol/Sample/ra
      -- 
    ra_7514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2707_inst_ack_0, ack => convTransposeD_CP_6792_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	1 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2701/phi_stmt_2701_sources/type_cast_2707/SplitProtocol/Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2701/phi_stmt_2701_sources/type_cast_2707/SplitProtocol/Update/ca
      -- 
    ca_7519_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2707_inst_ack_1, ack => convTransposeD_CP_6792_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	94 
    -- CP-element group 84:  members (5) 
      -- CP-element group 84: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2701/$exit
      -- CP-element group 84: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2701/phi_stmt_2701_sources/$exit
      -- CP-element group 84: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2701/phi_stmt_2701_sources/type_cast_2707/$exit
      -- CP-element group 84: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2701/phi_stmt_2701_sources/type_cast_2707/SplitProtocol/$exit
      -- CP-element group 84: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2701/phi_stmt_2701_req
      -- 
    phi_stmt_2701_req_7520_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2701_req_7520_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(84), ack => phi_stmt_2701_req_1); -- 
    convTransposeD_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(82) & convTransposeD_CP_6792_elements(83);
      gj_convTransposeD_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	1 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2708/phi_stmt_2708_sources/type_cast_2714/SplitProtocol/Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2708/phi_stmt_2708_sources/type_cast_2714/SplitProtocol/Sample/ra
      -- 
    ra_7537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2714_inst_ack_0, ack => convTransposeD_CP_6792_elements(85)); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	1 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2708/phi_stmt_2708_sources/type_cast_2714/SplitProtocol/Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2708/phi_stmt_2708_sources/type_cast_2714/SplitProtocol/Update/ca
      -- 
    ca_7542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2714_inst_ack_1, ack => convTransposeD_CP_6792_elements(86)); -- 
    -- CP-element group 87:  join  transition  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	94 
    -- CP-element group 87:  members (5) 
      -- CP-element group 87: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2708/$exit
      -- CP-element group 87: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2708/phi_stmt_2708_sources/$exit
      -- CP-element group 87: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2708/phi_stmt_2708_sources/type_cast_2714/$exit
      -- CP-element group 87: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2708/phi_stmt_2708_sources/type_cast_2714/SplitProtocol/$exit
      -- CP-element group 87: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2708/phi_stmt_2708_req
      -- 
    phi_stmt_2708_req_7543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2708_req_7543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(87), ack => phi_stmt_2708_req_1); -- 
    convTransposeD_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(85) & convTransposeD_CP_6792_elements(86);
      gj_convTransposeD_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	1 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2715/phi_stmt_2715_sources/type_cast_2721/SplitProtocol/Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2715/phi_stmt_2715_sources/type_cast_2721/SplitProtocol/Sample/ra
      -- 
    ra_7560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2721_inst_ack_0, ack => convTransposeD_CP_6792_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	1 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2715/phi_stmt_2715_sources/type_cast_2721/SplitProtocol/Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2715/phi_stmt_2715_sources/type_cast_2721/SplitProtocol/Update/ca
      -- 
    ca_7565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2721_inst_ack_1, ack => convTransposeD_CP_6792_elements(89)); -- 
    -- CP-element group 90:  join  transition  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	94 
    -- CP-element group 90:  members (5) 
      -- CP-element group 90: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2715/$exit
      -- CP-element group 90: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2715/phi_stmt_2715_sources/$exit
      -- CP-element group 90: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2715/phi_stmt_2715_sources/type_cast_2721/$exit
      -- CP-element group 90: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2715/phi_stmt_2715_sources/type_cast_2721/SplitProtocol/$exit
      -- CP-element group 90: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2715/phi_stmt_2715_req
      -- 
    phi_stmt_2715_req_7566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2715_req_7566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(90), ack => phi_stmt_2715_req_1); -- 
    convTransposeD_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(88) & convTransposeD_CP_6792_elements(89);
      gj_convTransposeD_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	1 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2722/phi_stmt_2722_sources/type_cast_2727/SplitProtocol/Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2722/phi_stmt_2722_sources/type_cast_2727/SplitProtocol/Sample/ra
      -- 
    ra_7583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2727_inst_ack_0, ack => convTransposeD_CP_6792_elements(91)); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	1 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2722/phi_stmt_2722_sources/type_cast_2727/SplitProtocol/Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2722/phi_stmt_2722_sources/type_cast_2727/SplitProtocol/Update/ca
      -- 
    ca_7588_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2727_inst_ack_1, ack => convTransposeD_CP_6792_elements(92)); -- 
    -- CP-element group 93:  join  transition  output  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (5) 
      -- CP-element group 93: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2722/$exit
      -- CP-element group 93: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2722/phi_stmt_2722_sources/$exit
      -- CP-element group 93: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2722/phi_stmt_2722_sources/type_cast_2727/$exit
      -- CP-element group 93: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2722/phi_stmt_2722_sources/type_cast_2727/SplitProtocol/$exit
      -- CP-element group 93: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2722/phi_stmt_2722_req
      -- 
    phi_stmt_2722_req_7589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2722_req_7589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(93), ack => phi_stmt_2722_req_1); -- 
    convTransposeD_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(91) & convTransposeD_CP_6792_elements(92);
      gj_convTransposeD_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  join  transition  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	84 
    -- CP-element group 94: 	87 
    -- CP-element group 94: 	90 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (1) 
      -- CP-element group 94: 	 branch_block_stmt_2585/ifx_xend132_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(84) & convTransposeD_CP_6792_elements(87) & convTransposeD_CP_6792_elements(90) & convTransposeD_CP_6792_elements(93);
      gj_convTransposeD_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  merge  fork  transition  place  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	81 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95: 	97 
    -- CP-element group 95: 	98 
    -- CP-element group 95: 	99 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_2585/merge_stmt_2700_PhiReqMerge
      -- CP-element group 95: 	 branch_block_stmt_2585/merge_stmt_2700_PhiAck/$entry
      -- 
    convTransposeD_CP_6792_elements(95) <= OrReduce(convTransposeD_CP_6792_elements(81) & convTransposeD_CP_6792_elements(94));
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	100 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_2585/merge_stmt_2700_PhiAck/phi_stmt_2701_ack
      -- 
    phi_stmt_2701_ack_7594_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2701_ack_0, ack => convTransposeD_CP_6792_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	100 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_2585/merge_stmt_2700_PhiAck/phi_stmt_2708_ack
      -- 
    phi_stmt_2708_ack_7595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2708_ack_0, ack => convTransposeD_CP_6792_elements(97)); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	95 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	100 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_2585/merge_stmt_2700_PhiAck/phi_stmt_2715_ack
      -- 
    phi_stmt_2715_ack_7596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2715_ack_0, ack => convTransposeD_CP_6792_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	95 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_2585/merge_stmt_2700_PhiAck/phi_stmt_2722_ack
      -- 
    phi_stmt_2722_ack_7597_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2722_ack_0, ack => convTransposeD_CP_6792_elements(99)); -- 
    -- CP-element group 100:  join  fork  transition  place  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	96 
    -- CP-element group 100: 	97 
    -- CP-element group 100: 	98 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	42 
    -- CP-element group 100: 	43 
    -- CP-element group 100: 	44 
    -- CP-element group 100: 	45 
    -- CP-element group 100: 	46 
    -- CP-element group 100: 	47 
    -- CP-element group 100: 	48 
    -- CP-element group 100: 	49 
    -- CP-element group 100: 	51 
    -- CP-element group 100: 	53 
    -- CP-element group 100: 	55 
    -- CP-element group 100: 	58 
    -- CP-element group 100: 	60 
    -- CP-element group 100: 	63 
    -- CP-element group 100: 	64 
    -- CP-element group 100: 	65 
    -- CP-element group 100:  members (56) 
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850__entry__
      -- CP-element group 100: 	 branch_block_stmt_2585/merge_stmt_2700__exit__
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2766_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2762_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2800_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2800_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2762_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2762_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2762_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2766_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/addr_of_2807_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/$entry
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2800_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2766_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2800_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2800_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2770_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2770_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2770_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2770_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2806_final_index_sum_regn_update_start
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/addr_of_2807_complete/$entry
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/addr_of_2807_complete/req
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2811_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2800_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2806_final_index_sum_regn_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2806_final_index_sum_regn_Update/req
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2766_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2766_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2770_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2770_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2766_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2762_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2762_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2811_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2811_Update/word_access_complete/$entry
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2811_Update/word_access_complete/word_0/$entry
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2811_Update/word_access_complete/word_0/cr
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/addr_of_2830_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2829_final_index_sum_regn_update_start
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2829_final_index_sum_regn_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/array_obj_ref_2829_final_index_sum_regn_Update/req
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/addr_of_2830_complete/$entry
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/addr_of_2830_complete/req
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2833_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2833_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2833_Update/word_access_complete/$entry
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2833_Update/word_access_complete/word_0/$entry
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/ptr_deref_2833_Update/word_access_complete/word_0/cr
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2838_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2838_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2838_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2838_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2838_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2585/assign_stmt_2734_to_assign_stmt_2850/type_cast_2838_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2585/merge_stmt_2700_PhiAck/$exit
      -- 
    rr_7154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(100), ack => type_cast_2800_inst_req_0); -- 
    cr_7117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(100), ack => type_cast_2762_inst_req_1); -- 
    cr_7159_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7159_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(100), ack => type_cast_2800_inst_req_1); -- 
    rr_7126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(100), ack => type_cast_2766_inst_req_0); -- 
    rr_7140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(100), ack => type_cast_2770_inst_req_0); -- 
    req_7205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(100), ack => addr_of_2807_final_reg_req_1); -- 
    req_7190_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7190_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(100), ack => array_obj_ref_2806_index_offset_req_1); -- 
    cr_7145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(100), ack => type_cast_2770_inst_req_1); -- 
    cr_7131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(100), ack => type_cast_2766_inst_req_1); -- 
    rr_7112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(100), ack => type_cast_2762_inst_req_0); -- 
    cr_7250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(100), ack => ptr_deref_2811_load_0_req_1); -- 
    req_7286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(100), ack => array_obj_ref_2829_index_offset_req_1); -- 
    req_7301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(100), ack => addr_of_2830_final_reg_req_1); -- 
    cr_7351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(100), ack => ptr_deref_2833_store_0_req_1); -- 
    rr_7360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(100), ack => type_cast_2838_inst_req_0); -- 
    cr_7365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(100), ack => type_cast_2838_inst_req_1); -- 
    convTransposeD_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(96) & convTransposeD_CP_6792_elements(97) & convTransposeD_CP_6792_elements(98) & convTransposeD_CP_6792_elements(99);
      gj_convTransposeD_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  transition  output  delay-element  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	72 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	108 
    -- CP-element group 101:  members (4) 
      -- CP-element group 101: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2905/$exit
      -- CP-element group 101: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2905/phi_stmt_2905_sources/$exit
      -- CP-element group 101: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2905/phi_stmt_2905_sources/type_cast_2911_konst_delay_trans
      -- CP-element group 101: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2905/phi_stmt_2905_req
      -- 
    phi_stmt_2905_req_7632_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2905_req_7632_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(101), ack => phi_stmt_2905_req_1); -- 
    -- Element group convTransposeD_CP_6792_elements(101) is a control-delay.
    cp_element_101_delay: control_delay_element  generic map(name => " 101_delay", delay_value => 1)  port map(req => convTransposeD_CP_6792_elements(72), ack => convTransposeD_CP_6792_elements(101), clk => clk, reset =>reset);
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	72 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2912/phi_stmt_2912_sources/type_cast_2917/SplitProtocol/Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2912/phi_stmt_2912_sources/type_cast_2917/SplitProtocol/Sample/ra
      -- 
    ra_7649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2917_inst_ack_0, ack => convTransposeD_CP_6792_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	72 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2912/phi_stmt_2912_sources/type_cast_2917/SplitProtocol/Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2912/phi_stmt_2912_sources/type_cast_2917/SplitProtocol/Update/ca
      -- 
    ca_7654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2917_inst_ack_1, ack => convTransposeD_CP_6792_elements(103)); -- 
    -- CP-element group 104:  join  transition  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	108 
    -- CP-element group 104:  members (5) 
      -- CP-element group 104: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2912/$exit
      -- CP-element group 104: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2912/phi_stmt_2912_sources/$exit
      -- CP-element group 104: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2912/phi_stmt_2912_sources/type_cast_2917/$exit
      -- CP-element group 104: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2912/phi_stmt_2912_sources/type_cast_2917/SplitProtocol/$exit
      -- CP-element group 104: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2912/phi_stmt_2912_req
      -- 
    phi_stmt_2912_req_7655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2912_req_7655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(104), ack => phi_stmt_2912_req_1); -- 
    convTransposeD_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(102) & convTransposeD_CP_6792_elements(103);
      gj_convTransposeD_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	72 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2923/SplitProtocol/Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2923/SplitProtocol/Sample/ra
      -- 
    ra_7672_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2923_inst_ack_0, ack => convTransposeD_CP_6792_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	72 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2923/SplitProtocol/Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2923/SplitProtocol/Update/ca
      -- 
    ca_7677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2923_inst_ack_1, ack => convTransposeD_CP_6792_elements(106)); -- 
    -- CP-element group 107:  join  transition  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (5) 
      -- CP-element group 107: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2918/$exit
      -- CP-element group 107: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/$exit
      -- CP-element group 107: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2923/$exit
      -- CP-element group 107: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2923/SplitProtocol/$exit
      -- CP-element group 107: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_req
      -- 
    phi_stmt_2918_req_7678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2918_req_7678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(107), ack => phi_stmt_2918_req_1); -- 
    convTransposeD_cp_element_group_107: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_107"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(105) & convTransposeD_CP_6792_elements(106);
      gj_convTransposeD_cp_element_group_107 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 108:  join  transition  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	101 
    -- CP-element group 108: 	104 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	119 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_2585/ifx_xelse_ifx_xend132_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(101) & convTransposeD_CP_6792_elements(104) & convTransposeD_CP_6792_elements(107);
      gj_convTransposeD_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	67 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2905/phi_stmt_2905_sources/type_cast_2908/SplitProtocol/Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2905/phi_stmt_2905_sources/type_cast_2908/SplitProtocol/Sample/ra
      -- 
    ra_7698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2908_inst_ack_0, ack => convTransposeD_CP_6792_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	67 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2905/phi_stmt_2905_sources/type_cast_2908/SplitProtocol/Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2905/phi_stmt_2905_sources/type_cast_2908/SplitProtocol/Update/ca
      -- 
    ca_7703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2908_inst_ack_1, ack => convTransposeD_CP_6792_elements(110)); -- 
    -- CP-element group 111:  join  transition  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	118 
    -- CP-element group 111:  members (5) 
      -- CP-element group 111: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2905/$exit
      -- CP-element group 111: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2905/phi_stmt_2905_sources/$exit
      -- CP-element group 111: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2905/phi_stmt_2905_sources/type_cast_2908/$exit
      -- CP-element group 111: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2905/phi_stmt_2905_sources/type_cast_2908/SplitProtocol/$exit
      -- CP-element group 111: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2905/phi_stmt_2905_req
      -- 
    phi_stmt_2905_req_7704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2905_req_7704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(111), ack => phi_stmt_2905_req_0); -- 
    convTransposeD_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(109) & convTransposeD_CP_6792_elements(110);
      gj_convTransposeD_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	67 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (2) 
      -- CP-element group 112: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2912/phi_stmt_2912_sources/type_cast_2915/SplitProtocol/Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2912/phi_stmt_2912_sources/type_cast_2915/SplitProtocol/Sample/ra
      -- 
    ra_7721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2915_inst_ack_0, ack => convTransposeD_CP_6792_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	67 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2912/phi_stmt_2912_sources/type_cast_2915/SplitProtocol/Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2912/phi_stmt_2912_sources/type_cast_2915/SplitProtocol/Update/ca
      -- 
    ca_7726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2915_inst_ack_1, ack => convTransposeD_CP_6792_elements(113)); -- 
    -- CP-element group 114:  join  transition  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	118 
    -- CP-element group 114:  members (5) 
      -- CP-element group 114: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2912/$exit
      -- CP-element group 114: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2912/phi_stmt_2912_sources/$exit
      -- CP-element group 114: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2912/phi_stmt_2912_sources/type_cast_2915/$exit
      -- CP-element group 114: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2912/phi_stmt_2912_sources/type_cast_2915/SplitProtocol/$exit
      -- CP-element group 114: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2912/phi_stmt_2912_req
      -- 
    phi_stmt_2912_req_7727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2912_req_7727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(114), ack => phi_stmt_2912_req_0); -- 
    convTransposeD_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(112) & convTransposeD_CP_6792_elements(113);
      gj_convTransposeD_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	67 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2921/SplitProtocol/Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2921/SplitProtocol/Sample/ra
      -- 
    ra_7744_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2921_inst_ack_0, ack => convTransposeD_CP_6792_elements(115)); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	67 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116:  members (2) 
      -- CP-element group 116: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2921/SplitProtocol/Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2921/SplitProtocol/Update/ca
      -- 
    ca_7749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2921_inst_ack_1, ack => convTransposeD_CP_6792_elements(116)); -- 
    -- CP-element group 117:  join  transition  output  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (5) 
      -- CP-element group 117: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2918/$exit
      -- CP-element group 117: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/$exit
      -- CP-element group 117: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2921/$exit
      -- CP-element group 117: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2921/SplitProtocol/$exit
      -- CP-element group 117: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_req
      -- 
    phi_stmt_2918_req_7750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2918_req_7750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(117), ack => phi_stmt_2918_req_0); -- 
    convTransposeD_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(115) & convTransposeD_CP_6792_elements(116);
      gj_convTransposeD_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  join  transition  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	111 
    -- CP-element group 118: 	114 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_2585/ifx_xthen_ifx_xend132_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(111) & convTransposeD_CP_6792_elements(114) & convTransposeD_CP_6792_elements(117);
      gj_convTransposeD_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  merge  fork  transition  place  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	108 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119: 	121 
    -- CP-element group 119: 	122 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_2585/merge_stmt_2904_PhiReqMerge
      -- CP-element group 119: 	 branch_block_stmt_2585/merge_stmt_2904_PhiAck/$entry
      -- 
    convTransposeD_CP_6792_elements(119) <= OrReduce(convTransposeD_CP_6792_elements(108) & convTransposeD_CP_6792_elements(118));
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	123 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_2585/merge_stmt_2904_PhiAck/phi_stmt_2905_ack
      -- 
    phi_stmt_2905_ack_7755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2905_ack_0, ack => convTransposeD_CP_6792_elements(120)); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	123 
    -- CP-element group 121:  members (1) 
      -- CP-element group 121: 	 branch_block_stmt_2585/merge_stmt_2904_PhiAck/phi_stmt_2912_ack
      -- 
    phi_stmt_2912_ack_7756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2912_ack_0, ack => convTransposeD_CP_6792_elements(121)); -- 
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	119 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_2585/merge_stmt_2904_PhiAck/phi_stmt_2918_ack
      -- 
    phi_stmt_2918_ack_7757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2918_ack_0, ack => convTransposeD_CP_6792_elements(122)); -- 
    -- CP-element group 123:  join  transition  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	120 
    -- CP-element group 123: 	121 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	1 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_2585/merge_stmt_2904_PhiAck/$exit
      -- 
    convTransposeD_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(120) & convTransposeD_CP_6792_elements(121) & convTransposeD_CP_6792_elements(122);
      gj_convTransposeD_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(123), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom91_2828_resized : std_logic_vector(13 downto 0);
    signal R_idxprom91_2828_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2805_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2805_scaled : std_logic_vector(13 downto 0);
    signal add103_2863 : std_logic_vector(15 downto 0);
    signal add32_2664 : std_logic_vector(15 downto 0);
    signal add50_2670 : std_logic_vector(15 downto 0);
    signal add63_2681 : std_logic_vector(15 downto 0);
    signal add82_2781 : std_logic_vector(63 downto 0);
    signal add84_2791 : std_logic_vector(63 downto 0);
    signal add96_2845 : std_logic_vector(31 downto 0);
    signal add_2637 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_2739 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2806_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2806_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2806_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2806_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2806_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2806_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2829_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2829_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2829_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2829_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2829_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2829_root_address : std_logic_vector(13 downto 0);
    signal arrayidx87_2808 : std_logic_vector(31 downto 0);
    signal arrayidx92_2831 : std_logic_vector(31 downto 0);
    signal call11_2606 : std_logic_vector(15 downto 0);
    signal call13_2609 : std_logic_vector(15 downto 0);
    signal call14_2612 : std_logic_vector(15 downto 0);
    signal call15_2615 : std_logic_vector(15 downto 0);
    signal call16_2628 : std_logic_vector(15 downto 0);
    signal call18_2640 : std_logic_vector(15 downto 0);
    signal call1_2591 : std_logic_vector(15 downto 0);
    signal call20_2643 : std_logic_vector(15 downto 0);
    signal call22_2646 : std_logic_vector(15 downto 0);
    signal call3_2594 : std_logic_vector(15 downto 0);
    signal call5_2597 : std_logic_vector(15 downto 0);
    signal call7_2600 : std_logic_vector(15 downto 0);
    signal call9_2603 : std_logic_vector(15 downto 0);
    signal call_2588 : std_logic_vector(15 downto 0);
    signal cmp111_2876 : std_logic_vector(0 downto 0);
    signal cmp121_2897 : std_logic_vector(0 downto 0);
    signal cmp_2850 : std_logic_vector(0 downto 0);
    signal conv17_2632 : std_logic_vector(31 downto 0);
    signal conv70_2763 : std_logic_vector(63 downto 0);
    signal conv73_2690 : std_logic_vector(63 downto 0);
    signal conv75_2767 : std_logic_vector(63 downto 0);
    signal conv78_2694 : std_logic_vector(63 downto 0);
    signal conv80_2771 : std_logic_vector(63 downto 0);
    signal conv95_2839 : std_logic_vector(31 downto 0);
    signal conv99_2698 : std_logic_vector(31 downto 0);
    signal conv_2619 : std_logic_vector(31 downto 0);
    signal idxprom91_2824 : std_logic_vector(63 downto 0);
    signal idxprom_2801 : std_logic_vector(63 downto 0);
    signal inc115_2880 : std_logic_vector(15 downto 0);
    signal inc115x_xinput_dim0x_x2_2885 : std_logic_vector(15 downto 0);
    signal inc_2871 : std_logic_vector(15 downto 0);
    signal indvar_2701 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_2930 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_2918 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_2722 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_2912 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_2715 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2892 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_2905 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2708 : std_logic_vector(15 downto 0);
    signal mul59_2754 : std_logic_vector(15 downto 0);
    signal mul81_2776 : std_logic_vector(63 downto 0);
    signal mul83_2786 : std_logic_vector(63 downto 0);
    signal mul_2744 : std_logic_vector(15 downto 0);
    signal ptr_deref_2811_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2811_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2811_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2811_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2811_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2833_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2833_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2833_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2833_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2833_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2833_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_2625 : std_logic_vector(31 downto 0);
    signal shr135_2653 : std_logic_vector(15 downto 0);
    signal shr31136_2659 : std_logic_vector(15 downto 0);
    signal shr86_2797 : std_logic_vector(31 downto 0);
    signal shr90_2818 : std_logic_vector(63 downto 0);
    signal sub53_2749 : std_logic_vector(15 downto 0);
    signal sub66_2686 : std_logic_vector(15 downto 0);
    signal sub67_2759 : std_logic_vector(15 downto 0);
    signal sub_2675 : std_logic_vector(15 downto 0);
    signal tmp1_2734 : std_logic_vector(31 downto 0);
    signal tmp88_2812 : std_logic_vector(63 downto 0);
    signal type_cast_2623_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2651_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2657_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2668_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2679_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2705_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2707_wire : std_logic_vector(31 downto 0);
    signal type_cast_2712_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2714_wire : std_logic_vector(15 downto 0);
    signal type_cast_2719_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2721_wire : std_logic_vector(15 downto 0);
    signal type_cast_2725_wire : std_logic_vector(15 downto 0);
    signal type_cast_2727_wire : std_logic_vector(15 downto 0);
    signal type_cast_2732_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2795_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2816_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2822_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2843_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2861_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2869_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2889_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2908_wire : std_logic_vector(15 downto 0);
    signal type_cast_2911_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2915_wire : std_logic_vector(15 downto 0);
    signal type_cast_2917_wire : std_logic_vector(15 downto 0);
    signal type_cast_2921_wire : std_logic_vector(15 downto 0);
    signal type_cast_2923_wire : std_logic_vector(15 downto 0);
    signal type_cast_2928_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2936_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_2806_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2806_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2806_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2806_resized_base_address <= "00000000000000";
    array_obj_ref_2829_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2829_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2829_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2829_resized_base_address <= "00000000000000";
    ptr_deref_2811_word_offset_0 <= "00000000000000";
    ptr_deref_2833_word_offset_0 <= "00000000000000";
    type_cast_2623_wire_constant <= "00000000000000000000000000010000";
    type_cast_2651_wire_constant <= "0000000000000010";
    type_cast_2657_wire_constant <= "0000000000000001";
    type_cast_2668_wire_constant <= "1111111111111111";
    type_cast_2679_wire_constant <= "1111111111111111";
    type_cast_2705_wire_constant <= "00000000000000000000000000000000";
    type_cast_2712_wire_constant <= "0000000000000000";
    type_cast_2719_wire_constant <= "0000000000000000";
    type_cast_2732_wire_constant <= "00000000000000000000000000000100";
    type_cast_2795_wire_constant <= "00000000000000000000000000000010";
    type_cast_2816_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_2822_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_2843_wire_constant <= "00000000000000000000000000000100";
    type_cast_2861_wire_constant <= "0000000000000100";
    type_cast_2869_wire_constant <= "0000000000000001";
    type_cast_2889_wire_constant <= "0000000000000000";
    type_cast_2911_wire_constant <= "0000000000000000";
    type_cast_2928_wire_constant <= "00000000000000000000000000000001";
    type_cast_2936_wire_constant <= "0000000000000001";
    phi_stmt_2701: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2705_wire_constant & type_cast_2707_wire;
      req <= phi_stmt_2701_req_0 & phi_stmt_2701_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2701",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2701_ack_0,
          idata => idata,
          odata => indvar_2701,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2701
    phi_stmt_2708: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2712_wire_constant & type_cast_2714_wire;
      req <= phi_stmt_2708_req_0 & phi_stmt_2708_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2708",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2708_ack_0,
          idata => idata,
          odata => input_dim2x_x1_2708,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2708
    phi_stmt_2715: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2719_wire_constant & type_cast_2721_wire;
      req <= phi_stmt_2715_req_0 & phi_stmt_2715_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2715",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2715_ack_0,
          idata => idata,
          odata => input_dim1x_x1_2715,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2715
    phi_stmt_2722: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2725_wire & type_cast_2727_wire;
      req <= phi_stmt_2722_req_0 & phi_stmt_2722_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2722",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2722_ack_0,
          idata => idata,
          odata => input_dim0x_x2_2722,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2722
    phi_stmt_2905: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2908_wire & type_cast_2911_wire_constant;
      req <= phi_stmt_2905_req_0 & phi_stmt_2905_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2905",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2905_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_2905,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2905
    phi_stmt_2912: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2915_wire & type_cast_2917_wire;
      req <= phi_stmt_2912_req_0 & phi_stmt_2912_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2912",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2912_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_2912,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2912
    phi_stmt_2918: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2921_wire & type_cast_2923_wire;
      req <= phi_stmt_2918_req_0 & phi_stmt_2918_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2918",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2918_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_2918,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2918
    -- flow-through select operator MUX_2891_inst
    input_dim1x_x2_2892 <= type_cast_2889_wire_constant when (cmp111_2876(0) /=  '0') else inc_2871;
    addr_of_2807_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2807_final_reg_req_0;
      addr_of_2807_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2807_final_reg_req_1;
      addr_of_2807_final_reg_ack_1<= rack(0);
      addr_of_2807_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2807_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2806_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx87_2808,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2830_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2830_final_reg_req_0;
      addr_of_2830_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2830_final_reg_req_1;
      addr_of_2830_final_reg_ack_1<= rack(0);
      addr_of_2830_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2830_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2829_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx92_2831,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2618_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2618_inst_req_0;
      type_cast_2618_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2618_inst_req_1;
      type_cast_2618_inst_ack_1<= rack(0);
      type_cast_2618_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2618_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_2615,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_2619,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2631_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2631_inst_req_0;
      type_cast_2631_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2631_inst_req_1;
      type_cast_2631_inst_ack_1<= rack(0);
      type_cast_2631_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2631_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_2628,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_2632,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2689_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2689_inst_req_0;
      type_cast_2689_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2689_inst_req_1;
      type_cast_2689_inst_ack_1<= rack(0);
      type_cast_2689_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2689_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_2646,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_2690,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2693_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2693_inst_req_0;
      type_cast_2693_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2693_inst_req_1;
      type_cast_2693_inst_ack_1<= rack(0);
      type_cast_2693_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2693_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_2643,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv78_2694,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2697_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2697_inst_req_0;
      type_cast_2697_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2697_inst_req_1;
      type_cast_2697_inst_ack_1<= rack(0);
      type_cast_2697_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2697_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_2594,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv99_2698,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2707_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2707_inst_req_0;
      type_cast_2707_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2707_inst_req_1;
      type_cast_2707_inst_ack_1<= rack(0);
      type_cast_2707_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2707_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2930,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2707_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2714_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2714_inst_req_0;
      type_cast_2714_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2714_inst_req_1;
      type_cast_2714_inst_ack_1<= rack(0);
      type_cast_2714_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2714_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_2905,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2714_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2721_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2721_inst_req_0;
      type_cast_2721_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2721_inst_req_1;
      type_cast_2721_inst_ack_1<= rack(0);
      type_cast_2721_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2721_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_2912,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2721_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2725_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2725_inst_req_0;
      type_cast_2725_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2725_inst_req_1;
      type_cast_2725_inst_ack_1<= rack(0);
      type_cast_2725_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2725_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add32_2664,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2725_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2727_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2727_inst_req_0;
      type_cast_2727_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2727_inst_req_1;
      type_cast_2727_inst_ack_1<= rack(0);
      type_cast_2727_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2727_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_2918,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2727_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2762_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2762_inst_req_0;
      type_cast_2762_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2762_inst_req_1;
      type_cast_2762_inst_ack_1<= rack(0);
      type_cast_2762_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2762_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2708,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_2763,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2766_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2766_inst_req_0;
      type_cast_2766_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2766_inst_req_1;
      type_cast_2766_inst_ack_1<= rack(0);
      type_cast_2766_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2766_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub67_2759,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_2767,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2770_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2770_inst_req_0;
      type_cast_2770_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2770_inst_req_1;
      type_cast_2770_inst_ack_1<= rack(0);
      type_cast_2770_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2770_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub53_2749,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv80_2771,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2800_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2800_inst_req_0;
      type_cast_2800_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2800_inst_req_1;
      type_cast_2800_inst_ack_1<= rack(0);
      type_cast_2800_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2800_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr86_2797,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2801,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2838_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2838_inst_req_0;
      type_cast_2838_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2838_inst_req_1;
      type_cast_2838_inst_ack_1<= rack(0);
      type_cast_2838_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2838_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2708,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_2839,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2879_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2879_inst_req_0;
      type_cast_2879_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2879_inst_req_1;
      type_cast_2879_inst_ack_1<= rack(0);
      type_cast_2879_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2879_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp111_2876,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc115_2880,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2908_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2908_inst_req_0;
      type_cast_2908_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2908_inst_req_1;
      type_cast_2908_inst_ack_1<= rack(0);
      type_cast_2908_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2908_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add103_2863,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2908_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2915_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2915_inst_req_0;
      type_cast_2915_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2915_inst_req_1;
      type_cast_2915_inst_ack_1<= rack(0);
      type_cast_2915_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2915_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_2715,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2915_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2917_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2917_inst_req_0;
      type_cast_2917_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2917_inst_req_1;
      type_cast_2917_inst_ack_1<= rack(0);
      type_cast_2917_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2917_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2892,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2917_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2921_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2921_inst_req_0;
      type_cast_2921_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2921_inst_req_1;
      type_cast_2921_inst_ack_1<= rack(0);
      type_cast_2921_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2921_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_2722,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2921_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2923_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2923_inst_req_0;
      type_cast_2923_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2923_inst_req_1;
      type_cast_2923_inst_ack_1<= rack(0);
      type_cast_2923_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2923_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc115x_xinput_dim0x_x2_2885,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2923_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_2806_index_1_rename
    process(R_idxprom_2805_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2805_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2805_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2806_index_1_resize
    process(idxprom_2801) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2801;
      ov := iv(13 downto 0);
      R_idxprom_2805_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2806_root_address_inst
    process(array_obj_ref_2806_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2806_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2806_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2829_index_1_rename
    process(R_idxprom91_2828_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom91_2828_resized;
      ov(13 downto 0) := iv;
      R_idxprom91_2828_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2829_index_1_resize
    process(idxprom91_2824) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom91_2824;
      ov := iv(13 downto 0);
      R_idxprom91_2828_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2829_root_address_inst
    process(array_obj_ref_2829_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2829_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2829_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2811_addr_0
    process(ptr_deref_2811_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2811_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2811_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2811_base_resize
    process(arrayidx87_2808) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx87_2808;
      ov := iv(13 downto 0);
      ptr_deref_2811_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2811_gather_scatter
    process(ptr_deref_2811_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2811_data_0;
      ov(63 downto 0) := iv;
      tmp88_2812 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2811_root_address_inst
    process(ptr_deref_2811_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2811_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2811_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2833_addr_0
    process(ptr_deref_2833_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2833_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2833_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2833_base_resize
    process(arrayidx92_2831) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx92_2831;
      ov := iv(13 downto 0);
      ptr_deref_2833_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2833_gather_scatter
    process(tmp88_2812) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp88_2812;
      ov(63 downto 0) := iv;
      ptr_deref_2833_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2833_root_address_inst
    process(ptr_deref_2833_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2833_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2833_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2851_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2850;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2851_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2851_branch_req_0,
          ack0 => if_stmt_2851_branch_ack_0,
          ack1 => if_stmt_2851_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2898_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp121_2897;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2898_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2898_branch_req_0,
          ack0 => if_stmt_2898_branch_ack_0,
          ack1 => if_stmt_2898_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2663_inst
    process(shr135_2653, shr31136_2659) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr135_2653, shr31136_2659, tmp_var);
      add32_2664 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2669_inst
    process(call7_2600) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_2600, type_cast_2668_wire_constant, tmp_var);
      add50_2670 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2680_inst
    process(call9_2603) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_2603, type_cast_2679_wire_constant, tmp_var);
      add63_2681 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2748_inst
    process(sub_2675, mul_2744) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_2675, mul_2744, tmp_var);
      sub53_2749 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2758_inst
    process(sub66_2686, mul59_2754) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub66_2686, mul59_2754, tmp_var);
      sub67_2759 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2862_inst
    process(input_dim2x_x1_2708) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_2708, type_cast_2861_wire_constant, tmp_var);
      add103_2863 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2870_inst
    process(input_dim1x_x1_2715) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_2715, type_cast_2869_wire_constant, tmp_var);
      inc_2871 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2884_inst
    process(inc115_2880, input_dim0x_x2_2722) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc115_2880, input_dim0x_x2_2722, tmp_var);
      inc115x_xinput_dim0x_x2_2885 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2738_inst
    process(add_2637, tmp1_2734) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_2637, tmp1_2734, tmp_var);
      add_src_0x_x0_2739 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2844_inst
    process(conv95_2839) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv95_2839, type_cast_2843_wire_constant, tmp_var);
      add96_2845 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2929_inst
    process(indvar_2701) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2701, type_cast_2928_wire_constant, tmp_var);
      indvarx_xnext_2930 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2780_inst
    process(mul81_2776, conv75_2767) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul81_2776, conv75_2767, tmp_var);
      add82_2781 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2790_inst
    process(mul83_2786, conv70_2763) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul83_2786, conv70_2763, tmp_var);
      add84_2791 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2823_inst
    process(shr90_2818) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr90_2818, type_cast_2822_wire_constant, tmp_var);
      idxprom91_2824 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2875_inst
    process(inc_2871, call1_2591) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_2871, call1_2591, tmp_var);
      cmp111_2876 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2896_inst
    process(inc115x_xinput_dim0x_x2_2885, call_2588) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc115x_xinput_dim0x_x2_2885, call_2588, tmp_var);
      cmp121_2897 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2652_inst
    process(call_2588) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_2588, type_cast_2651_wire_constant, tmp_var);
      shr135_2653 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2658_inst
    process(call_2588) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_2588, type_cast_2657_wire_constant, tmp_var);
      shr31136_2659 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2796_inst
    process(add_src_0x_x0_2739) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_2739, type_cast_2795_wire_constant, tmp_var);
      shr86_2797 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2817_inst
    process(add84_2791) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add84_2791, type_cast_2816_wire_constant, tmp_var);
      shr90_2818 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2743_inst
    process(input_dim0x_x2_2722, call13_2609) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x2_2722, call13_2609, tmp_var);
      mul_2744 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2753_inst
    process(input_dim1x_x1_2715, call13_2609) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_2715, call13_2609, tmp_var);
      mul59_2754 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2733_inst
    process(indvar_2701) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2701, type_cast_2732_wire_constant, tmp_var);
      tmp1_2734 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2775_inst
    process(conv80_2771, conv78_2694) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv80_2771, conv78_2694, tmp_var);
      mul81_2776 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2785_inst
    process(add82_2781, conv73_2690) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add82_2781, conv73_2690, tmp_var);
      mul83_2786 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_2636_inst
    process(shl_2625, conv17_2632) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_2625, conv17_2632, tmp_var);
      add_2637 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2624_inst
    process(conv_2619) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_2619, type_cast_2623_wire_constant, tmp_var);
      shl_2625 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2674_inst
    process(add50_2670, call14_2612) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add50_2670, call14_2612, tmp_var);
      sub_2675 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2685_inst
    process(add63_2681, call14_2612) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add63_2681, call14_2612, tmp_var);
      sub66_2686 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2849_inst
    process(add96_2845, conv99_2698) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add96_2845, conv99_2698, tmp_var);
      cmp_2850 <= tmp_var; --
    end process;
    -- shared split operator group (30) : array_obj_ref_2806_index_offset 
    ApIntAdd_group_30: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2805_scaled;
      array_obj_ref_2806_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2806_index_offset_req_0;
      array_obj_ref_2806_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2806_index_offset_req_1;
      array_obj_ref_2806_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_30_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_30_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_30",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared split operator group (31) : array_obj_ref_2829_index_offset 
    ApIntAdd_group_31: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom91_2828_scaled;
      array_obj_ref_2829_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2829_index_offset_req_0;
      array_obj_ref_2829_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2829_index_offset_req_1;
      array_obj_ref_2829_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_31_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_31_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_31",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared load operator group (0) : ptr_deref_2811_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2811_load_0_req_0;
      ptr_deref_2811_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2811_load_0_req_1;
      ptr_deref_2811_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2811_word_address_0;
      ptr_deref_2811_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_2833_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2833_store_0_req_0;
      ptr_deref_2833_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2833_store_0_req_1;
      ptr_deref_2833_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2833_word_address_0;
      data_in <= ptr_deref_2833_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block3_start_2587_inst RPIPE_Block3_start_2590_inst RPIPE_Block3_start_2593_inst RPIPE_Block3_start_2596_inst RPIPE_Block3_start_2599_inst RPIPE_Block3_start_2602_inst RPIPE_Block3_start_2605_inst RPIPE_Block3_start_2608_inst RPIPE_Block3_start_2611_inst RPIPE_Block3_start_2614_inst RPIPE_Block3_start_2627_inst RPIPE_Block3_start_2639_inst RPIPE_Block3_start_2642_inst RPIPE_Block3_start_2645_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block3_start_2587_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block3_start_2590_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block3_start_2593_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block3_start_2596_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block3_start_2599_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block3_start_2602_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block3_start_2605_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block3_start_2608_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block3_start_2611_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block3_start_2614_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block3_start_2627_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block3_start_2639_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block3_start_2642_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block3_start_2645_inst_req_0;
      RPIPE_Block3_start_2587_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block3_start_2590_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block3_start_2593_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block3_start_2596_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block3_start_2599_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block3_start_2602_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block3_start_2605_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block3_start_2608_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block3_start_2611_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block3_start_2614_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block3_start_2627_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block3_start_2639_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block3_start_2642_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block3_start_2645_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block3_start_2587_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block3_start_2590_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block3_start_2593_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block3_start_2596_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block3_start_2599_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block3_start_2602_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block3_start_2605_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block3_start_2608_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block3_start_2611_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block3_start_2614_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block3_start_2627_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block3_start_2639_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block3_start_2642_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block3_start_2645_inst_req_1;
      RPIPE_Block3_start_2587_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block3_start_2590_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block3_start_2593_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block3_start_2596_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block3_start_2599_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block3_start_2602_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block3_start_2605_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block3_start_2608_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block3_start_2611_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block3_start_2614_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block3_start_2627_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block3_start_2639_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block3_start_2642_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block3_start_2645_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call_2588 <= data_out(223 downto 208);
      call1_2591 <= data_out(207 downto 192);
      call3_2594 <= data_out(191 downto 176);
      call5_2597 <= data_out(175 downto 160);
      call7_2600 <= data_out(159 downto 144);
      call9_2603 <= data_out(143 downto 128);
      call11_2606 <= data_out(127 downto 112);
      call13_2609 <= data_out(111 downto 96);
      call14_2612 <= data_out(95 downto 80);
      call15_2615 <= data_out(79 downto 64);
      call16_2628 <= data_out(63 downto 48);
      call18_2640 <= data_out(47 downto 32);
      call20_2643 <= data_out(31 downto 16);
      call22_2646 <= data_out(15 downto 0);
      Block3_start_read_0_gI: SplitGuardInterface generic map(name => "Block3_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_start_read_0: InputPortRevised -- 
        generic map ( name => "Block3_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_start_pipe_read_req(0),
          oack => Block3_start_pipe_read_ack(0),
          odata => Block3_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block3_done_2934_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block3_done_2934_inst_req_0;
      WPIPE_Block3_done_2934_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block3_done_2934_inst_req_1;
      WPIPE_Block3_done_2934_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2936_wire_constant;
      Block3_done_write_0_gI: SplitGuardInterface generic map(name => "Block3_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block3_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_done_pipe_write_req(0),
          oack => Block3_done_pipe_write_ack(0),
          odata => Block3_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeD_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    c : out  std_logic_vector(63 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal c_buffer :  std_logic_vector(63 downto 0);
  signal c_update_enable: Boolean;
  signal timer_CP_0_start: Boolean;
  signal timer_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal LOAD_count_29_load_0_req_0 : boolean;
  signal LOAD_count_29_load_0_ack_0 : boolean;
  signal LOAD_count_29_load_0_req_1 : boolean;
  signal LOAD_count_29_load_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= c_buffer;
  c <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_0: Block -- control-path 
    signal timer_CP_0_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    timer_CP_0_elements(0) <= timer_CP_0_start;
    timer_CP_0_symbol <= timer_CP_0_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_Update/$entry
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_30/$entry
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_sample_start_
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_update_start_
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_Sample/$entry
      -- 
    rr_21_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_21_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => LOAD_count_29_load_0_req_0); -- 
    cr_32_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_32_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => LOAD_count_29_load_0_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 assign_stmt_30/LOAD_count_29_Sample/word_access_start/$exit
      -- CP-element group 1: 	 assign_stmt_30/LOAD_count_29_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 assign_stmt_30/LOAD_count_29_Sample/word_access_start/word_0/ra
      -- CP-element group 1: 	 assign_stmt_30/LOAD_count_29_sample_completed_
      -- CP-element group 1: 	 assign_stmt_30/LOAD_count_29_Sample/$exit
      -- 
    ra_22_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_29_load_0_ack_0, ack => timer_CP_0_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_Update/$exit
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_Update/word_access_complete/$exit
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_Update/LOAD_count_29_Merge/$entry
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_30/$exit
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_update_completed_
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_Update/LOAD_count_29_Merge/$exit
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_Update/LOAD_count_29_Merge/merge_req
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_Update/LOAD_count_29_Merge/merge_ack
      -- 
    ca_33_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_29_load_0_ack_1, ack => timer_CP_0_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_count_29_data_0 : std_logic_vector(63 downto 0);
    signal LOAD_count_29_word_address_0 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    LOAD_count_29_word_address_0 <= "0";
    -- equivalence LOAD_count_29_gather_scatter
    process(LOAD_count_29_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_count_29_data_0;
      ov(63 downto 0) := iv;
      c_buffer <= ov(63 downto 0);
      --
    end process;
    -- shared load operator group (0) : LOAD_count_29_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_count_29_load_0_req_0;
      LOAD_count_29_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_count_29_load_0_req_1;
      LOAD_count_29_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_count_29_word_address_0;
      LOAD_count_29_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(0 downto 0),
          mtag => memory_space_0_lr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    ConvTranspose_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    ConvTranspose_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    ConvTranspose_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_read_data: out std_logic_vector(63 downto 0);
    elapsed_time_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(55 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(75 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(255 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(10 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_3
  signal memory_space_3_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_3_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_3_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_3_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_3_sr_req :  std_logic_vector(4 downto 0);
  signal memory_space_3_sr_ack : std_logic_vector(4 downto 0);
  signal memory_space_3_sr_addr : std_logic_vector(69 downto 0);
  signal memory_space_3_sr_data : std_logic_vector(319 downto 0);
  signal memory_space_3_sr_tag : std_logic_vector(94 downto 0);
  signal memory_space_3_sc_req : std_logic_vector(4 downto 0);
  signal memory_space_3_sc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_3_sc_tag :  std_logic_vector(4 downto 0);
  -- declarations related to module convTranspose
  component convTranspose is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTranspose
  signal convTranspose_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTranspose_tag_out   : std_logic_vector(1 downto 0);
  signal convTranspose_start_req : std_logic;
  signal convTranspose_start_ack : std_logic;
  signal convTranspose_fin_req   : std_logic;
  signal convTranspose_fin_ack : std_logic;
  -- declarations related to module convTransposeA
  component convTransposeA is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeA
  signal convTransposeA_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeA_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeA_start_req : std_logic;
  signal convTransposeA_start_ack : std_logic;
  signal convTransposeA_fin_req   : std_logic;
  signal convTransposeA_fin_ack : std_logic;
  -- declarations related to module convTransposeB
  component convTransposeB is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeB
  signal convTransposeB_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeB_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeB_start_req : std_logic;
  signal convTransposeB_start_ack : std_logic;
  signal convTransposeB_fin_req   : std_logic;
  signal convTransposeB_fin_ack : std_logic;
  -- declarations related to module convTransposeC
  component convTransposeC is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeC
  signal convTransposeC_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeC_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeC_start_req : std_logic;
  signal convTransposeC_start_ack : std_logic;
  signal convTransposeC_fin_req   : std_logic;
  signal convTransposeC_fin_ack : std_logic;
  -- declarations related to module convTransposeD
  component convTransposeD is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeD
  signal convTransposeD_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeD_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeD_start_req : std_logic;
  signal convTransposeD_start_ack : std_logic;
  signal convTransposeD_fin_req   : std_logic;
  signal convTransposeD_fin_ack : std_logic;
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_c :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe Block0_done
  signal Block0_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_done
  signal Block0_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block0_start
  signal Block0_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_start
  signal Block0_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_done
  signal Block1_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_done
  signal Block1_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_start
  signal Block1_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_start
  signal Block1_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_done
  signal Block2_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_done
  signal Block2_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_start
  signal Block2_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_start
  signal Block2_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_done
  signal Block3_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_done
  signal Block3_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_start
  signal Block3_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_start
  signal Block3_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe ConvTranspose_input_pipe
  signal ConvTranspose_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe ConvTranspose_output_pipe
  signal ConvTranspose_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe elapsed_time_pipe
  signal elapsed_time_pipe_pipe_write_data: std_logic_vector(63 downto 0);
  signal elapsed_time_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal elapsed_time_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module convTranspose
  convTranspose_instance:convTranspose-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTranspose_start_req,
      start_ack => convTranspose_start_ack,
      fin_req => convTranspose_fin_req,
      fin_ack => convTranspose_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_3_lr_req => memory_space_3_lr_req(0 downto 0),
      memory_space_3_lr_ack => memory_space_3_lr_ack(0 downto 0),
      memory_space_3_lr_addr => memory_space_3_lr_addr(13 downto 0),
      memory_space_3_lr_tag => memory_space_3_lr_tag(18 downto 0),
      memory_space_3_lc_req => memory_space_3_lc_req(0 downto 0),
      memory_space_3_lc_ack => memory_space_3_lc_ack(0 downto 0),
      memory_space_3_lc_data => memory_space_3_lc_data(63 downto 0),
      memory_space_3_lc_tag => memory_space_3_lc_tag(0 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(18 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(0 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(10 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(63 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(0 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(0 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(4 downto 4),
      memory_space_3_sr_ack => memory_space_3_sr_ack(4 downto 4),
      memory_space_3_sr_addr => memory_space_3_sr_addr(69 downto 56),
      memory_space_3_sr_data => memory_space_3_sr_data(319 downto 256),
      memory_space_3_sr_tag => memory_space_3_sr_tag(94 downto 76),
      memory_space_3_sc_req => memory_space_3_sc_req(4 downto 4),
      memory_space_3_sc_ack => memory_space_3_sc_ack(4 downto 4),
      memory_space_3_sc_tag => memory_space_3_sc_tag(4 downto 4),
      Block0_done_pipe_read_req => Block0_done_pipe_read_req(0 downto 0),
      Block0_done_pipe_read_ack => Block0_done_pipe_read_ack(0 downto 0),
      Block0_done_pipe_read_data => Block0_done_pipe_read_data(15 downto 0),
      Block1_done_pipe_read_req => Block1_done_pipe_read_req(0 downto 0),
      Block1_done_pipe_read_ack => Block1_done_pipe_read_ack(0 downto 0),
      Block1_done_pipe_read_data => Block1_done_pipe_read_data(15 downto 0),
      ConvTranspose_input_pipe_pipe_read_req => ConvTranspose_input_pipe_pipe_read_req(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_ack => ConvTranspose_input_pipe_pipe_read_ack(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_data => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
      Block2_done_pipe_read_req => Block2_done_pipe_read_req(0 downto 0),
      Block2_done_pipe_read_ack => Block2_done_pipe_read_ack(0 downto 0),
      Block2_done_pipe_read_data => Block2_done_pipe_read_data(15 downto 0),
      Block3_done_pipe_read_req => Block3_done_pipe_read_req(0 downto 0),
      Block3_done_pipe_read_ack => Block3_done_pipe_read_ack(0 downto 0),
      Block3_done_pipe_read_data => Block3_done_pipe_read_data(15 downto 0),
      Block1_start_pipe_write_req => Block1_start_pipe_write_req(0 downto 0),
      Block1_start_pipe_write_ack => Block1_start_pipe_write_ack(0 downto 0),
      Block1_start_pipe_write_data => Block1_start_pipe_write_data(15 downto 0),
      Block0_start_pipe_write_req => Block0_start_pipe_write_req(0 downto 0),
      Block0_start_pipe_write_ack => Block0_start_pipe_write_ack(0 downto 0),
      Block0_start_pipe_write_data => Block0_start_pipe_write_data(15 downto 0),
      Block3_start_pipe_write_req => Block3_start_pipe_write_req(0 downto 0),
      Block3_start_pipe_write_ack => Block3_start_pipe_write_ack(0 downto 0),
      Block3_start_pipe_write_data => Block3_start_pipe_write_data(15 downto 0),
      ConvTranspose_output_pipe_pipe_write_req => ConvTranspose_output_pipe_pipe_write_req(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_ack => ConvTranspose_output_pipe_pipe_write_ack(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_data => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
      Block2_start_pipe_write_req => Block2_start_pipe_write_req(0 downto 0),
      Block2_start_pipe_write_ack => Block2_start_pipe_write_ack(0 downto 0),
      Block2_start_pipe_write_data => Block2_start_pipe_write_data(15 downto 0),
      elapsed_time_pipe_pipe_write_req => elapsed_time_pipe_pipe_write_req(0 downto 0),
      elapsed_time_pipe_pipe_write_ack => elapsed_time_pipe_pipe_write_ack(0 downto 0),
      elapsed_time_pipe_pipe_write_data => elapsed_time_pipe_pipe_write_data(63 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      tag_in => convTranspose_tag_in,
      tag_out => convTranspose_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTranspose_tag_in <= (others => '0');
  convTranspose_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTranspose_start_req, start_ack => convTranspose_start_ack,  fin_req => convTranspose_fin_req,  fin_ack => convTranspose_fin_ack);
  -- module convTransposeA
  convTransposeA_instance:convTransposeA-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeA_start_req,
      start_ack => convTransposeA_start_ack,
      fin_req => convTransposeA_fin_req,
      fin_ack => convTransposeA_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(3 downto 3),
      memory_space_1_lr_ack => memory_space_1_lr_ack(3 downto 3),
      memory_space_1_lr_addr => memory_space_1_lr_addr(55 downto 42),
      memory_space_1_lr_tag => memory_space_1_lr_tag(75 downto 57),
      memory_space_1_lc_req => memory_space_1_lc_req(3 downto 3),
      memory_space_1_lc_ack => memory_space_1_lc_ack(3 downto 3),
      memory_space_1_lc_data => memory_space_1_lc_data(255 downto 192),
      memory_space_1_lc_tag => memory_space_1_lc_tag(3 downto 3),
      memory_space_3_sr_req => memory_space_3_sr_req(3 downto 3),
      memory_space_3_sr_ack => memory_space_3_sr_ack(3 downto 3),
      memory_space_3_sr_addr => memory_space_3_sr_addr(55 downto 42),
      memory_space_3_sr_data => memory_space_3_sr_data(255 downto 192),
      memory_space_3_sr_tag => memory_space_3_sr_tag(75 downto 57),
      memory_space_3_sc_req => memory_space_3_sc_req(3 downto 3),
      memory_space_3_sc_ack => memory_space_3_sc_ack(3 downto 3),
      memory_space_3_sc_tag => memory_space_3_sc_tag(3 downto 3),
      Block0_start_pipe_read_req => Block0_start_pipe_read_req(0 downto 0),
      Block0_start_pipe_read_ack => Block0_start_pipe_read_ack(0 downto 0),
      Block0_start_pipe_read_data => Block0_start_pipe_read_data(15 downto 0),
      Block0_done_pipe_write_req => Block0_done_pipe_write_req(0 downto 0),
      Block0_done_pipe_write_ack => Block0_done_pipe_write_ack(0 downto 0),
      Block0_done_pipe_write_data => Block0_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeA_tag_in,
      tag_out => convTransposeA_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeA_tag_in <= (others => '0');
  convTransposeA_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeA_start_req, start_ack => convTransposeA_start_ack,  fin_req => convTransposeA_fin_req,  fin_ack => convTransposeA_fin_ack);
  -- module convTransposeB
  convTransposeB_instance:convTransposeB-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeB_start_req,
      start_ack => convTransposeB_start_ack,
      fin_req => convTransposeB_fin_req,
      fin_ack => convTransposeB_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(2 downto 2),
      memory_space_1_lr_ack => memory_space_1_lr_ack(2 downto 2),
      memory_space_1_lr_addr => memory_space_1_lr_addr(41 downto 28),
      memory_space_1_lr_tag => memory_space_1_lr_tag(56 downto 38),
      memory_space_1_lc_req => memory_space_1_lc_req(2 downto 2),
      memory_space_1_lc_ack => memory_space_1_lc_ack(2 downto 2),
      memory_space_1_lc_data => memory_space_1_lc_data(191 downto 128),
      memory_space_1_lc_tag => memory_space_1_lc_tag(2 downto 2),
      memory_space_3_sr_req => memory_space_3_sr_req(2 downto 2),
      memory_space_3_sr_ack => memory_space_3_sr_ack(2 downto 2),
      memory_space_3_sr_addr => memory_space_3_sr_addr(41 downto 28),
      memory_space_3_sr_data => memory_space_3_sr_data(191 downto 128),
      memory_space_3_sr_tag => memory_space_3_sr_tag(56 downto 38),
      memory_space_3_sc_req => memory_space_3_sc_req(2 downto 2),
      memory_space_3_sc_ack => memory_space_3_sc_ack(2 downto 2),
      memory_space_3_sc_tag => memory_space_3_sc_tag(2 downto 2),
      Block1_start_pipe_read_req => Block1_start_pipe_read_req(0 downto 0),
      Block1_start_pipe_read_ack => Block1_start_pipe_read_ack(0 downto 0),
      Block1_start_pipe_read_data => Block1_start_pipe_read_data(15 downto 0),
      Block1_done_pipe_write_req => Block1_done_pipe_write_req(0 downto 0),
      Block1_done_pipe_write_ack => Block1_done_pipe_write_ack(0 downto 0),
      Block1_done_pipe_write_data => Block1_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeB_tag_in,
      tag_out => convTransposeB_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeB_tag_in <= (others => '0');
  convTransposeB_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeB_start_req, start_ack => convTransposeB_start_ack,  fin_req => convTransposeB_fin_req,  fin_ack => convTransposeB_fin_ack);
  -- module convTransposeC
  convTransposeC_instance:convTransposeC-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeC_start_req,
      start_ack => convTransposeC_start_ack,
      fin_req => convTransposeC_fin_req,
      fin_ack => convTransposeC_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(1 downto 1),
      memory_space_1_lr_ack => memory_space_1_lr_ack(1 downto 1),
      memory_space_1_lr_addr => memory_space_1_lr_addr(27 downto 14),
      memory_space_1_lr_tag => memory_space_1_lr_tag(37 downto 19),
      memory_space_1_lc_req => memory_space_1_lc_req(1 downto 1),
      memory_space_1_lc_ack => memory_space_1_lc_ack(1 downto 1),
      memory_space_1_lc_data => memory_space_1_lc_data(127 downto 64),
      memory_space_1_lc_tag => memory_space_1_lc_tag(1 downto 1),
      memory_space_3_sr_req => memory_space_3_sr_req(1 downto 1),
      memory_space_3_sr_ack => memory_space_3_sr_ack(1 downto 1),
      memory_space_3_sr_addr => memory_space_3_sr_addr(27 downto 14),
      memory_space_3_sr_data => memory_space_3_sr_data(127 downto 64),
      memory_space_3_sr_tag => memory_space_3_sr_tag(37 downto 19),
      memory_space_3_sc_req => memory_space_3_sc_req(1 downto 1),
      memory_space_3_sc_ack => memory_space_3_sc_ack(1 downto 1),
      memory_space_3_sc_tag => memory_space_3_sc_tag(1 downto 1),
      Block2_start_pipe_read_req => Block2_start_pipe_read_req(0 downto 0),
      Block2_start_pipe_read_ack => Block2_start_pipe_read_ack(0 downto 0),
      Block2_start_pipe_read_data => Block2_start_pipe_read_data(15 downto 0),
      Block2_done_pipe_write_req => Block2_done_pipe_write_req(0 downto 0),
      Block2_done_pipe_write_ack => Block2_done_pipe_write_ack(0 downto 0),
      Block2_done_pipe_write_data => Block2_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeC_tag_in,
      tag_out => convTransposeC_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeC_tag_in <= (others => '0');
  convTransposeC_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeC_start_req, start_ack => convTransposeC_start_ack,  fin_req => convTransposeC_fin_req,  fin_ack => convTransposeC_fin_ack);
  -- module convTransposeD
  convTransposeD_instance:convTransposeD-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeD_start_req,
      start_ack => convTransposeD_start_ack,
      fin_req => convTransposeD_fin_req,
      fin_ack => convTransposeD_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(18 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(0 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(0 downto 0),
      memory_space_3_sr_ack => memory_space_3_sr_ack(0 downto 0),
      memory_space_3_sr_addr => memory_space_3_sr_addr(13 downto 0),
      memory_space_3_sr_data => memory_space_3_sr_data(63 downto 0),
      memory_space_3_sr_tag => memory_space_3_sr_tag(18 downto 0),
      memory_space_3_sc_req => memory_space_3_sc_req(0 downto 0),
      memory_space_3_sc_ack => memory_space_3_sc_ack(0 downto 0),
      memory_space_3_sc_tag => memory_space_3_sc_tag(0 downto 0),
      Block3_start_pipe_read_req => Block3_start_pipe_read_req(0 downto 0),
      Block3_start_pipe_read_ack => Block3_start_pipe_read_ack(0 downto 0),
      Block3_start_pipe_read_data => Block3_start_pipe_read_data(15 downto 0),
      Block3_done_pipe_write_req => Block3_done_pipe_write_req(0 downto 0),
      Block3_done_pipe_write_ack => Block3_done_pipe_write_ack(0 downto 0),
      Block3_done_pipe_write_data => Block3_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeD_tag_in,
      tag_out => convTransposeD_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeD_tag_in <= (others => '0');
  convTransposeD_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeD_start_req, start_ack => convTransposeD_start_ack,  fin_req => convTransposeD_fin_req,  fin_ack => convTransposeD_fin_ack);
  -- module timer
  timer_out_args <= timer_c ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      c => timer_c,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(0 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(0 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  Block0_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_done_pipe_read_req,
      read_ack => Block0_done_pipe_read_ack,
      read_data => Block0_done_pipe_read_data,
      write_req => Block0_done_pipe_write_req,
      write_ack => Block0_done_pipe_write_ack,
      write_data => Block0_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block0_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_start_pipe_read_req,
      read_ack => Block0_start_pipe_read_ack,
      read_data => Block0_start_pipe_read_data,
      write_req => Block0_start_pipe_write_req,
      write_ack => Block0_start_pipe_write_ack,
      write_data => Block0_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_done_pipe_read_req,
      read_ack => Block1_done_pipe_read_ack,
      read_data => Block1_done_pipe_read_data,
      write_req => Block1_done_pipe_write_req,
      write_ack => Block1_done_pipe_write_ack,
      write_data => Block1_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_start_pipe_read_req,
      read_ack => Block1_start_pipe_read_ack,
      read_data => Block1_start_pipe_read_data,
      write_req => Block1_start_pipe_write_req,
      write_ack => Block1_start_pipe_write_ack,
      write_data => Block1_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_done_pipe_read_req,
      read_ack => Block2_done_pipe_read_ack,
      read_data => Block2_done_pipe_read_data,
      write_req => Block2_done_pipe_write_req,
      write_ack => Block2_done_pipe_write_ack,
      write_data => Block2_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_start_pipe_read_req,
      read_ack => Block2_start_pipe_read_ack,
      read_data => Block2_start_pipe_read_data,
      write_req => Block2_start_pipe_write_req,
      write_ack => Block2_start_pipe_write_ack,
      write_data => Block2_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_done_pipe_read_req,
      read_ack => Block3_done_pipe_read_ack,
      read_data => Block3_done_pipe_read_data,
      write_req => Block3_done_pipe_write_req,
      write_ack => Block3_done_pipe_write_ack,
      write_data => Block3_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_start_pipe_read_req,
      read_ack => Block3_start_pipe_read_ack,
      read_data => Block3_start_pipe_read_data,
      write_req => Block3_start_pipe_write_req,
      write_ack => Block3_start_pipe_write_ack,
      write_data => Block3_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_input_pipe_pipe_read_req,
      read_ack => ConvTranspose_input_pipe_pipe_read_ack,
      read_data => ConvTranspose_input_pipe_pipe_read_data,
      write_req => ConvTranspose_input_pipe_pipe_write_req,
      write_ack => ConvTranspose_input_pipe_pipe_write_ack,
      write_data => ConvTranspose_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_output_pipe_pipe_read_req,
      read_ack => ConvTranspose_output_pipe_pipe_read_ack,
      read_data => ConvTranspose_output_pipe_pipe_read_data,
      write_req => ConvTranspose_output_pipe_pipe_write_req,
      write_ack => ConvTranspose_output_pipe_pipe_write_ack,
      write_data => ConvTranspose_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  elapsed_time_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe elapsed_time_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => elapsed_time_pipe_pipe_read_req,
      read_ack => elapsed_time_pipe_pipe_read_ack,
      read_data => elapsed_time_pipe_pipe_read_data,
      write_req => elapsed_time_pipe_pipe_write_req,
      write_ack => elapsed_time_pipe_pipe_write_ack,
      write_data => elapsed_time_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  dummyROM_memory_space_0: dummy_read_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      addr_width => 1,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 4,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_2: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_stores => 1,
      addr_width => 11,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_3: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_3",
      num_loads => 1,
      num_stores => 5,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_3_lr_addr,
      lr_req_in => memory_space_3_lr_req,
      lr_ack_out => memory_space_3_lr_ack,
      lr_tag_in => memory_space_3_lr_tag,
      lc_req_in => memory_space_3_lc_req,
      lc_ack_out => memory_space_3_lc_ack,
      lc_data_out => memory_space_3_lc_data,
      lc_tag_out => memory_space_3_lc_tag,
      sr_addr_in => memory_space_3_sr_addr,
      sr_data_in => memory_space_3_sr_data,
      sr_req_in => memory_space_3_sr_req,
      sr_ack_out => memory_space_3_sr_ack,
      sr_tag_in => memory_space_3_sr_tag,
      sc_req_in=> memory_space_3_sc_req,
      sc_ack_out => memory_space_3_sc_ack,
      sc_tag_out => memory_space_3_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
