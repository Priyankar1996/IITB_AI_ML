-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTranspose is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(10 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTranspose;
architecture convTranspose_arch of convTranspose is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTranspose_CP_39_start: Boolean;
  signal convTranspose_CP_39_symbol: Boolean;
  -- volatile/operator module components. 
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal WPIPE_ConvTranspose_output_pipe_1103_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_718_inst_req_1 : boolean;
  signal type_cast_1060_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_718_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_988_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_718_inst_req_0 : boolean;
  signal type_cast_1060_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_718_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_953_inst_req_1 : boolean;
  signal addr_of_666_final_reg_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1097_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1091_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_41_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_41_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_529_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_529_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_565_inst_ack_1 : boolean;
  signal type_cast_569_inst_ack_1 : boolean;
  signal type_cast_569_inst_req_1 : boolean;
  signal type_cast_515_inst_ack_1 : boolean;
  signal type_cast_515_inst_req_1 : boolean;
  signal type_cast_569_inst_ack_0 : boolean;
  signal type_cast_515_inst_ack_0 : boolean;
  signal type_cast_569_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_28_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_28_inst_ack_0 : boolean;
  signal if_stmt_609_branch_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_28_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_28_inst_ack_1 : boolean;
  signal type_cast_686_inst_req_1 : boolean;
  signal type_cast_32_inst_req_0 : boolean;
  signal type_cast_32_inst_ack_0 : boolean;
  signal type_cast_32_inst_req_1 : boolean;
  signal type_cast_32_inst_ack_1 : boolean;
  signal type_cast_704_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1097_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_41_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_41_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_959_inst_req_1 : boolean;
  signal WPIPE_Block0_start_950_inst_ack_1 : boolean;
  signal type_cast_132_inst_req_0 : boolean;
  signal type_cast_132_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1091_inst_req_0 : boolean;
  signal type_cast_132_inst_req_1 : boolean;
  signal type_cast_132_inst_ack_1 : boolean;
  signal type_cast_45_inst_req_0 : boolean;
  signal WPIPE_Block0_start_962_inst_req_0 : boolean;
  signal type_cast_45_inst_ack_0 : boolean;
  signal type_cast_45_inst_req_1 : boolean;
  signal type_cast_45_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_669_inst_ack_1 : boolean;
  signal type_cast_704_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_565_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_53_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_53_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_53_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_53_inst_ack_1 : boolean;
  signal type_cast_1060_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1094_inst_req_0 : boolean;
  signal WPIPE_Block0_start_950_inst_req_1 : boolean;
  signal RPIPE_Block0_done_993_inst_req_0 : boolean;
  signal type_cast_57_inst_req_0 : boolean;
  signal type_cast_57_inst_ack_0 : boolean;
  signal type_cast_57_inst_req_1 : boolean;
  signal type_cast_57_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_66_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_66_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_565_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_66_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_66_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_700_inst_ack_1 : boolean;
  signal if_stmt_609_branch_ack_1 : boolean;
  signal type_cast_70_inst_req_0 : boolean;
  signal type_cast_70_inst_ack_0 : boolean;
  signal type_cast_70_inst_req_1 : boolean;
  signal type_cast_70_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_669_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_565_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_78_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_78_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_78_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_78_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1103_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_682_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_968_inst_req_0 : boolean;
  signal type_cast_82_inst_req_0 : boolean;
  signal type_cast_82_inst_ack_0 : boolean;
  signal type_cast_82_inst_req_1 : boolean;
  signal type_cast_82_inst_ack_1 : boolean;
  signal type_cast_704_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_91_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_91_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_91_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_91_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_682_inst_req_1 : boolean;
  signal type_cast_686_inst_ack_0 : boolean;
  signal type_cast_95_inst_req_0 : boolean;
  signal type_cast_95_inst_ack_0 : boolean;
  signal type_cast_95_inst_req_1 : boolean;
  signal ptr_deref_595_store_0_ack_1 : boolean;
  signal type_cast_95_inst_ack_1 : boolean;
  signal type_cast_704_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_103_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_103_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_103_inst_req_1 : boolean;
  signal ptr_deref_595_store_0_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_103_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_700_inst_req_1 : boolean;
  signal WPIPE_Block0_start_965_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_682_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1094_inst_ack_0 : boolean;
  signal type_cast_686_inst_req_0 : boolean;
  signal RPIPE_Block0_done_993_inst_ack_0 : boolean;
  signal if_stmt_609_branch_req_0 : boolean;
  signal type_cast_107_inst_req_0 : boolean;
  signal type_cast_107_inst_ack_0 : boolean;
  signal type_cast_107_inst_req_1 : boolean;
  signal type_cast_107_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_669_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_116_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_116_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_116_inst_req_1 : boolean;
  signal WPIPE_Block0_start_968_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_116_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_682_inst_req_0 : boolean;
  signal type_cast_120_inst_req_0 : boolean;
  signal type_cast_120_inst_ack_0 : boolean;
  signal type_cast_120_inst_req_1 : boolean;
  signal type_cast_120_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_669_inst_req_0 : boolean;
  signal WPIPE_Block0_start_968_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_128_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_128_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_128_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_128_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_319_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_319_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1100_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_319_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_319_inst_ack_1 : boolean;
  signal call_stmt_997_call_req_0 : boolean;
  signal type_cast_323_inst_req_0 : boolean;
  signal type_cast_323_inst_ack_0 : boolean;
  signal type_cast_551_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_953_inst_req_0 : boolean;
  signal type_cast_636_inst_ack_1 : boolean;
  signal type_cast_636_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_141_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_141_inst_ack_0 : boolean;
  signal type_cast_551_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_141_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_141_inst_ack_1 : boolean;
  signal type_cast_587_inst_ack_1 : boolean;
  signal array_obj_ref_665_index_offset_ack_1 : boolean;
  signal type_cast_145_inst_req_0 : boolean;
  signal ptr_deref_595_store_0_ack_0 : boolean;
  signal type_cast_145_inst_ack_0 : boolean;
  signal type_cast_145_inst_req_1 : boolean;
  signal type_cast_145_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_988_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_153_inst_req_0 : boolean;
  signal ptr_deref_595_store_0_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_153_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_153_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_153_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_700_inst_ack_0 : boolean;
  signal array_obj_ref_665_index_offset_req_1 : boolean;
  signal type_cast_157_inst_req_0 : boolean;
  signal type_cast_157_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1091_inst_ack_1 : boolean;
  signal type_cast_157_inst_req_1 : boolean;
  signal type_cast_157_inst_ack_1 : boolean;
  signal type_cast_686_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_965_inst_req_1 : boolean;
  signal type_cast_551_inst_ack_0 : boolean;
  signal type_cast_636_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_166_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_166_inst_ack_0 : boolean;
  signal type_cast_551_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_166_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_166_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_968_inst_ack_1 : boolean;
  signal type_cast_587_inst_req_1 : boolean;
  signal type_cast_636_inst_req_0 : boolean;
  signal type_cast_170_inst_req_0 : boolean;
  signal type_cast_170_inst_ack_0 : boolean;
  signal type_cast_170_inst_req_1 : boolean;
  signal type_cast_170_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_953_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_178_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_178_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_178_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_178_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_700_inst_req_0 : boolean;
  signal RPIPE_Block0_done_993_inst_req_1 : boolean;
  signal RPIPE_Block0_done_993_inst_ack_1 : boolean;
  signal type_cast_587_inst_ack_0 : boolean;
  signal type_cast_182_inst_req_0 : boolean;
  signal type_cast_182_inst_ack_0 : boolean;
  signal array_obj_ref_665_index_offset_ack_0 : boolean;
  signal type_cast_182_inst_req_1 : boolean;
  signal type_cast_182_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_191_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_191_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_191_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_191_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_959_inst_ack_1 : boolean;
  signal addr_of_666_final_reg_ack_1 : boolean;
  signal type_cast_1060_inst_ack_1 : boolean;
  signal type_cast_587_inst_req_0 : boolean;
  signal type_cast_195_inst_req_0 : boolean;
  signal type_cast_195_inst_ack_0 : boolean;
  signal array_obj_ref_665_index_offset_req_0 : boolean;
  signal type_cast_195_inst_req_1 : boolean;
  signal type_cast_195_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_547_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_547_inst_req_1 : boolean;
  signal type_cast_204_inst_req_0 : boolean;
  signal type_cast_204_inst_ack_0 : boolean;
  signal type_cast_204_inst_req_1 : boolean;
  signal type_cast_204_inst_ack_1 : boolean;
  signal type_cast_208_inst_req_0 : boolean;
  signal type_cast_208_inst_ack_0 : boolean;
  signal type_cast_208_inst_req_1 : boolean;
  signal type_cast_208_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_547_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_547_inst_req_0 : boolean;
  signal type_cast_212_inst_req_0 : boolean;
  signal type_cast_212_inst_ack_0 : boolean;
  signal type_cast_212_inst_req_1 : boolean;
  signal type_cast_212_inst_ack_1 : boolean;
  signal type_cast_226_inst_req_0 : boolean;
  signal type_cast_226_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_511_inst_ack_1 : boolean;
  signal type_cast_226_inst_req_1 : boolean;
  signal type_cast_226_inst_ack_1 : boolean;
  signal type_cast_230_inst_req_0 : boolean;
  signal type_cast_230_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_511_inst_req_1 : boolean;
  signal type_cast_230_inst_req_1 : boolean;
  signal type_cast_230_inst_ack_1 : boolean;
  signal type_cast_234_inst_req_0 : boolean;
  signal type_cast_234_inst_ack_0 : boolean;
  signal type_cast_234_inst_req_1 : boolean;
  signal type_cast_234_inst_ack_1 : boolean;
  signal type_cast_533_inst_ack_1 : boolean;
  signal type_cast_533_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_583_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_583_inst_req_1 : boolean;
  signal type_cast_238_inst_req_0 : boolean;
  signal type_cast_238_inst_ack_0 : boolean;
  signal type_cast_238_inst_req_1 : boolean;
  signal type_cast_238_inst_ack_1 : boolean;
  signal type_cast_533_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_256_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_256_inst_ack_0 : boolean;
  signal type_cast_533_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_256_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_256_inst_ack_1 : boolean;
  signal type_cast_673_inst_ack_1 : boolean;
  signal type_cast_673_inst_req_1 : boolean;
  signal addr_of_666_final_reg_req_1 : boolean;
  signal type_cast_260_inst_req_0 : boolean;
  signal type_cast_260_inst_ack_0 : boolean;
  signal type_cast_260_inst_req_1 : boolean;
  signal type_cast_260_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_269_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_269_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_269_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_269_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_583_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_583_inst_req_0 : boolean;
  signal type_cast_273_inst_req_0 : boolean;
  signal type_cast_273_inst_ack_0 : boolean;
  signal type_cast_273_inst_req_1 : boolean;
  signal type_cast_273_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_281_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_281_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_281_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_281_inst_ack_1 : boolean;
  signal type_cast_673_inst_ack_0 : boolean;
  signal type_cast_285_inst_req_0 : boolean;
  signal type_cast_285_inst_ack_0 : boolean;
  signal type_cast_285_inst_req_1 : boolean;
  signal type_cast_285_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_529_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1091_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_529_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_294_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_294_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_294_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_294_inst_ack_1 : boolean;
  signal type_cast_673_inst_req_0 : boolean;
  signal addr_of_666_final_reg_ack_0 : boolean;
  signal type_cast_515_inst_req_0 : boolean;
  signal type_cast_298_inst_req_0 : boolean;
  signal type_cast_298_inst_ack_0 : boolean;
  signal type_cast_298_inst_req_1 : boolean;
  signal type_cast_298_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_306_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_306_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_306_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_306_inst_ack_1 : boolean;
  signal type_cast_310_inst_req_0 : boolean;
  signal type_cast_310_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_953_inst_ack_1 : boolean;
  signal type_cast_310_inst_req_1 : boolean;
  signal type_cast_310_inst_ack_1 : boolean;
  signal type_cast_323_inst_req_1 : boolean;
  signal type_cast_323_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_978_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1085_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_331_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_331_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_331_inst_req_1 : boolean;
  signal call_stmt_997_call_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_331_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1094_inst_req_1 : boolean;
  signal type_cast_335_inst_req_0 : boolean;
  signal type_cast_335_inst_ack_0 : boolean;
  signal type_cast_335_inst_req_1 : boolean;
  signal type_cast_335_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_971_inst_req_0 : boolean;
  signal WPIPE_Block0_start_971_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_344_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_344_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_344_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_344_inst_ack_1 : boolean;
  signal type_cast_348_inst_req_0 : boolean;
  signal type_cast_348_inst_ack_0 : boolean;
  signal type_cast_348_inst_req_1 : boolean;
  signal call_stmt_997_call_req_1 : boolean;
  signal type_cast_348_inst_ack_1 : boolean;
  signal type_cast_1020_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_356_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_356_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_356_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_356_inst_ack_1 : boolean;
  signal type_cast_360_inst_req_0 : boolean;
  signal type_cast_360_inst_ack_0 : boolean;
  signal type_cast_360_inst_req_1 : boolean;
  signal type_cast_360_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_971_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1085_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_369_inst_req_0 : boolean;
  signal type_cast_1070_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_369_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_369_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_369_inst_ack_1 : boolean;
  signal type_cast_1020_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_971_inst_ack_1 : boolean;
  signal call_stmt_997_call_ack_1 : boolean;
  signal type_cast_373_inst_req_0 : boolean;
  signal type_cast_1070_inst_ack_0 : boolean;
  signal type_cast_373_inst_ack_0 : boolean;
  signal type_cast_373_inst_req_1 : boolean;
  signal type_cast_373_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_978_inst_ack_0 : boolean;
  signal if_stmt_387_branch_req_0 : boolean;
  signal if_stmt_387_branch_ack_1 : boolean;
  signal if_stmt_387_branch_ack_0 : boolean;
  signal if_stmt_402_branch_req_0 : boolean;
  signal if_stmt_402_branch_ack_1 : boolean;
  signal if_stmt_402_branch_ack_0 : boolean;
  signal type_cast_429_inst_req_0 : boolean;
  signal type_cast_429_inst_ack_0 : boolean;
  signal type_cast_429_inst_req_1 : boolean;
  signal type_cast_429_inst_ack_1 : boolean;
  signal array_obj_ref_458_index_offset_req_0 : boolean;
  signal array_obj_ref_458_index_offset_ack_0 : boolean;
  signal array_obj_ref_458_index_offset_req_1 : boolean;
  signal array_obj_ref_458_index_offset_ack_1 : boolean;
  signal addr_of_459_final_reg_req_0 : boolean;
  signal addr_of_459_final_reg_ack_0 : boolean;
  signal addr_of_459_final_reg_req_1 : boolean;
  signal addr_of_459_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_462_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_462_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_462_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_462_inst_ack_1 : boolean;
  signal type_cast_466_inst_req_0 : boolean;
  signal type_cast_466_inst_ack_0 : boolean;
  signal type_cast_466_inst_req_1 : boolean;
  signal type_cast_466_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_475_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_475_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_475_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_475_inst_ack_1 : boolean;
  signal type_cast_479_inst_req_0 : boolean;
  signal type_cast_479_inst_ack_0 : boolean;
  signal type_cast_479_inst_req_1 : boolean;
  signal type_cast_479_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_493_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_493_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_493_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_493_inst_ack_1 : boolean;
  signal type_cast_497_inst_req_0 : boolean;
  signal type_cast_497_inst_ack_0 : boolean;
  signal type_cast_497_inst_req_1 : boolean;
  signal type_cast_497_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_511_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_511_inst_ack_0 : boolean;
  signal type_cast_722_inst_req_0 : boolean;
  signal type_cast_722_inst_ack_0 : boolean;
  signal type_cast_722_inst_req_1 : boolean;
  signal type_cast_722_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_965_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_736_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_736_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_965_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_736_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_736_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_988_inst_ack_0 : boolean;
  signal type_cast_1080_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_988_inst_req_0 : boolean;
  signal type_cast_740_inst_req_0 : boolean;
  signal type_cast_740_inst_ack_0 : boolean;
  signal type_cast_740_inst_req_1 : boolean;
  signal type_cast_740_inst_ack_1 : boolean;
  signal if_stmt_1107_branch_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_754_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_754_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_754_inst_req_1 : boolean;
  signal type_cast_1050_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_754_inst_ack_1 : boolean;
  signal type_cast_1080_inst_req_1 : boolean;
  signal type_cast_758_inst_req_0 : boolean;
  signal type_cast_1050_inst_req_1 : boolean;
  signal type_cast_758_inst_ack_0 : boolean;
  signal type_cast_758_inst_req_1 : boolean;
  signal type_cast_758_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1082_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_772_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_772_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_772_inst_req_1 : boolean;
  signal type_cast_1050_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_772_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1100_inst_ack_1 : boolean;
  signal type_cast_776_inst_req_0 : boolean;
  signal type_cast_1050_inst_req_0 : boolean;
  signal type_cast_776_inst_ack_0 : boolean;
  signal type_cast_776_inst_req_1 : boolean;
  signal type_cast_776_inst_ack_1 : boolean;
  signal type_cast_1080_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1082_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_790_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_790_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_790_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_790_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1100_inst_req_1 : boolean;
  signal type_cast_794_inst_req_0 : boolean;
  signal type_cast_794_inst_ack_0 : boolean;
  signal type_cast_794_inst_req_1 : boolean;
  signal type_cast_794_inst_ack_1 : boolean;
  signal if_stmt_1107_branch_ack_1 : boolean;
  signal type_cast_1080_inst_req_0 : boolean;
  signal type_cast_1040_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_985_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_985_inst_req_1 : boolean;
  signal WPIPE_Block0_start_974_inst_ack_1 : boolean;
  signal type_cast_1040_inst_req_1 : boolean;
  signal WPIPE_Block0_start_974_inst_req_1 : boolean;
  signal ptr_deref_802_store_0_req_0 : boolean;
  signal ptr_deref_802_store_0_ack_0 : boolean;
  signal WPIPE_Block0_start_959_inst_ack_0 : boolean;
  signal ptr_deref_802_store_0_req_1 : boolean;
  signal ptr_deref_802_store_0_ack_1 : boolean;
  signal WPIPE_Block0_start_985_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_985_inst_req_0 : boolean;
  signal WPIPE_Block0_start_959_inst_req_0 : boolean;
  signal if_stmt_816_branch_req_0 : boolean;
  signal type_cast_1010_inst_ack_1 : boolean;
  signal if_stmt_816_branch_ack_1 : boolean;
  signal type_cast_1010_inst_req_1 : boolean;
  signal if_stmt_816_branch_ack_0 : boolean;
  signal type_cast_827_inst_req_0 : boolean;
  signal type_cast_827_inst_ack_0 : boolean;
  signal type_cast_827_inst_req_1 : boolean;
  signal type_cast_1040_inst_ack_0 : boolean;
  signal type_cast_827_inst_ack_1 : boolean;
  signal type_cast_831_inst_req_0 : boolean;
  signal type_cast_831_inst_ack_0 : boolean;
  signal type_cast_1010_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1088_inst_ack_1 : boolean;
  signal type_cast_831_inst_req_1 : boolean;
  signal type_cast_1040_inst_req_0 : boolean;
  signal type_cast_831_inst_ack_1 : boolean;
  signal type_cast_835_inst_req_0 : boolean;
  signal type_cast_835_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1088_inst_req_1 : boolean;
  signal type_cast_835_inst_req_1 : boolean;
  signal type_cast_835_inst_ack_1 : boolean;
  signal type_cast_1010_inst_req_0 : boolean;
  signal if_stmt_853_branch_req_0 : boolean;
  signal if_stmt_853_branch_ack_1 : boolean;
  signal WPIPE_Block0_start_956_inst_ack_1 : boolean;
  signal if_stmt_853_branch_ack_0 : boolean;
  signal WPIPE_Block0_start_974_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1085_inst_ack_1 : boolean;
  signal type_cast_880_inst_req_0 : boolean;
  signal type_cast_880_inst_ack_0 : boolean;
  signal type_cast_880_inst_req_1 : boolean;
  signal type_cast_880_inst_ack_1 : boolean;
  signal if_stmt_1107_branch_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1085_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1082_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_956_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1103_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_982_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_982_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1103_inst_req_0 : boolean;
  signal type_cast_1001_inst_ack_1 : boolean;
  signal array_obj_ref_909_index_offset_req_0 : boolean;
  signal array_obj_ref_909_index_offset_ack_0 : boolean;
  signal WPIPE_Block0_start_962_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1097_inst_ack_1 : boolean;
  signal array_obj_ref_909_index_offset_req_1 : boolean;
  signal array_obj_ref_909_index_offset_ack_1 : boolean;
  signal type_cast_1030_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_962_inst_req_1 : boolean;
  signal type_cast_1030_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1088_inst_ack_0 : boolean;
  signal addr_of_910_final_reg_req_0 : boolean;
  signal addr_of_910_final_reg_ack_0 : boolean;
  signal addr_of_910_final_reg_req_1 : boolean;
  signal addr_of_910_final_reg_ack_1 : boolean;
  signal WPIPE_Block0_start_982_inst_ack_0 : boolean;
  signal type_cast_1030_inst_ack_0 : boolean;
  signal type_cast_1070_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1097_inst_req_1 : boolean;
  signal type_cast_1030_inst_req_0 : boolean;
  signal WPIPE_Block0_start_982_inst_req_0 : boolean;
  signal type_cast_1001_inst_req_1 : boolean;
  signal WPIPE_Block0_start_974_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1082_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1088_inst_req_0 : boolean;
  signal ptr_deref_913_store_0_req_0 : boolean;
  signal ptr_deref_913_store_0_ack_0 : boolean;
  signal ptr_deref_913_store_0_req_1 : boolean;
  signal ptr_deref_913_store_0_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1100_inst_ack_0 : boolean;
  signal if_stmt_928_branch_req_0 : boolean;
  signal WPIPE_Block0_start_956_inst_ack_0 : boolean;
  signal if_stmt_928_branch_ack_1 : boolean;
  signal type_cast_1001_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_956_inst_req_0 : boolean;
  signal if_stmt_928_branch_ack_0 : boolean;
  signal type_cast_1001_inst_req_0 : boolean;
  signal call_stmt_939_call_req_0 : boolean;
  signal call_stmt_939_call_ack_0 : boolean;
  signal call_stmt_939_call_req_1 : boolean;
  signal call_stmt_939_call_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1094_inst_ack_1 : boolean;
  signal type_cast_1070_inst_req_1 : boolean;
  signal WPIPE_Block0_start_978_inst_ack_1 : boolean;
  signal type_cast_944_inst_req_0 : boolean;
  signal type_cast_1020_inst_ack_1 : boolean;
  signal type_cast_944_inst_ack_0 : boolean;
  signal type_cast_944_inst_req_1 : boolean;
  signal type_cast_1020_inst_req_1 : boolean;
  signal type_cast_944_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_978_inst_req_1 : boolean;
  signal WPIPE_Block0_start_950_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_947_inst_req_0 : boolean;
  signal WPIPE_Block0_start_947_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_962_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_947_inst_req_1 : boolean;
  signal WPIPE_Block0_start_947_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_950_inst_req_0 : boolean;
  signal type_cast_1134_inst_req_0 : boolean;
  signal type_cast_1134_inst_ack_0 : boolean;
  signal type_cast_1134_inst_req_1 : boolean;
  signal type_cast_1134_inst_ack_1 : boolean;
  signal array_obj_ref_1163_index_offset_req_0 : boolean;
  signal array_obj_ref_1163_index_offset_ack_0 : boolean;
  signal array_obj_ref_1163_index_offset_req_1 : boolean;
  signal array_obj_ref_1163_index_offset_ack_1 : boolean;
  signal addr_of_1164_final_reg_req_0 : boolean;
  signal addr_of_1164_final_reg_ack_0 : boolean;
  signal addr_of_1164_final_reg_req_1 : boolean;
  signal addr_of_1164_final_reg_ack_1 : boolean;
  signal ptr_deref_1168_load_0_req_0 : boolean;
  signal ptr_deref_1168_load_0_ack_0 : boolean;
  signal ptr_deref_1168_load_0_req_1 : boolean;
  signal ptr_deref_1168_load_0_ack_1 : boolean;
  signal phi_stmt_1151_ack_0 : boolean;
  signal type_cast_1172_inst_req_0 : boolean;
  signal type_cast_1172_inst_ack_0 : boolean;
  signal type_cast_1172_inst_req_1 : boolean;
  signal type_cast_1172_inst_ack_1 : boolean;
  signal type_cast_1182_inst_req_0 : boolean;
  signal type_cast_1182_inst_ack_0 : boolean;
  signal type_cast_1182_inst_req_1 : boolean;
  signal type_cast_1182_inst_ack_1 : boolean;
  signal type_cast_1192_inst_req_0 : boolean;
  signal type_cast_1192_inst_ack_0 : boolean;
  signal type_cast_1192_inst_req_1 : boolean;
  signal type_cast_1192_inst_ack_1 : boolean;
  signal type_cast_1202_inst_req_0 : boolean;
  signal type_cast_1202_inst_ack_0 : boolean;
  signal type_cast_1202_inst_req_1 : boolean;
  signal type_cast_1202_inst_ack_1 : boolean;
  signal type_cast_1212_inst_req_0 : boolean;
  signal type_cast_1212_inst_ack_0 : boolean;
  signal type_cast_1212_inst_req_1 : boolean;
  signal type_cast_1212_inst_ack_1 : boolean;
  signal type_cast_1222_inst_req_0 : boolean;
  signal type_cast_1222_inst_ack_0 : boolean;
  signal type_cast_1222_inst_req_1 : boolean;
  signal type_cast_1222_inst_ack_1 : boolean;
  signal type_cast_1232_inst_req_0 : boolean;
  signal type_cast_1232_inst_ack_0 : boolean;
  signal type_cast_1232_inst_req_1 : boolean;
  signal type_cast_1232_inst_ack_1 : boolean;
  signal type_cast_1242_inst_req_0 : boolean;
  signal type_cast_1242_inst_ack_0 : boolean;
  signal type_cast_1242_inst_req_1 : boolean;
  signal type_cast_1242_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1244_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1244_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1244_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1244_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1247_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1247_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1247_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1247_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1250_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1250_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1250_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1250_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1253_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1253_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1253_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1253_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1256_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1256_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1256_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1256_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1259_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1259_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1259_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1259_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1262_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1262_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1262_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1262_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1265_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1265_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1265_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1265_inst_ack_1 : boolean;
  signal if_stmt_1279_branch_req_0 : boolean;
  signal if_stmt_1279_branch_ack_1 : boolean;
  signal if_stmt_1279_branch_ack_0 : boolean;
  signal phi_stmt_446_req_0 : boolean;
  signal type_cast_452_inst_req_0 : boolean;
  signal type_cast_452_inst_ack_0 : boolean;
  signal type_cast_452_inst_req_1 : boolean;
  signal type_cast_452_inst_ack_1 : boolean;
  signal phi_stmt_446_req_1 : boolean;
  signal phi_stmt_446_ack_0 : boolean;
  signal phi_stmt_653_req_0 : boolean;
  signal type_cast_659_inst_req_0 : boolean;
  signal type_cast_659_inst_ack_0 : boolean;
  signal type_cast_659_inst_req_1 : boolean;
  signal type_cast_659_inst_ack_1 : boolean;
  signal phi_stmt_653_req_1 : boolean;
  signal phi_stmt_653_ack_0 : boolean;
  signal phi_stmt_897_req_0 : boolean;
  signal type_cast_903_inst_req_0 : boolean;
  signal type_cast_903_inst_ack_0 : boolean;
  signal type_cast_903_inst_req_1 : boolean;
  signal type_cast_903_inst_ack_1 : boolean;
  signal phi_stmt_897_req_1 : boolean;
  signal phi_stmt_897_ack_0 : boolean;
  signal phi_stmt_1151_req_0 : boolean;
  signal type_cast_1157_inst_req_0 : boolean;
  signal type_cast_1157_inst_ack_0 : boolean;
  signal type_cast_1157_inst_req_1 : boolean;
  signal type_cast_1157_inst_ack_1 : boolean;
  signal phi_stmt_1151_req_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTranspose_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTranspose_CP_39_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTranspose_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_39_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTranspose_CP_39_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_39_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTranspose_CP_39: Block -- control-path 
    signal convTranspose_CP_39_elements: BooleanArray(387 downto 0);
    -- 
  begin -- 
    convTranspose_CP_39_elements(0) <= convTranspose_CP_39_start;
    convTranspose_CP_39_symbol <= convTranspose_CP_39_elements(387);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	56 
    -- CP-element group 0: 	59 
    -- CP-element group 0: 	62 
    -- CP-element group 0: 	44 
    -- CP-element group 0: 	48 
    -- CP-element group 0: 	52 
    -- CP-element group 0: 	40 
    -- CP-element group 0: 	65 
    -- CP-element group 0: 	68 
    -- CP-element group 0: 	71 
    -- CP-element group 0: 	74 
    -- CP-element group 0: 	77 
    -- CP-element group 0: 	81 
    -- CP-element group 0: 	85 
    -- CP-element group 0: 	89 
    -- CP-element group 0: 	93 
    -- CP-element group 0: 	97 
    -- CP-element group 0: 	101 
    -- CP-element group 0: 	105 
    -- CP-element group 0: 	109 
    -- CP-element group 0: 	113 
    -- CP-element group 0: 	117 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	12 
    -- CP-element group 0: 	16 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	24 
    -- CP-element group 0: 	28 
    -- CP-element group 0: 	32 
    -- CP-element group 0: 	36 
    -- CP-element group 0:  members (101) 
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_26/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/branch_block_stmt_26__entry__
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_28_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_28_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_28_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_32_update_start_
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_32_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_32_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_132_update_start_
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_132_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_132_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_45_update_start_
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_45_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_45_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_57_update_start_
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_57_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_57_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_70_update_start_
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_70_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_70_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_82_update_start_
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_82_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_82_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_95_update_start_
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_95_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_95_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_107_update_start_
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_107_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_107_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_120_update_start_
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_120_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_120_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_323_update_start_
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_323_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_145_update_start_
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_145_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_145_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_157_update_start_
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_298_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_157_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_157_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_170_update_start_
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_170_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_170_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_182_update_start_
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_182_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_182_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_195_update_start_
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_195_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_195_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_204_update_start_
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_204_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_204_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_208_update_start_
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_208_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_208_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_212_update_start_
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_212_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_212_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_226_update_start_
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_226_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_226_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_230_update_start_
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_230_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_230_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_234_update_start_
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_234_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_234_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_238_update_start_
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_238_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_238_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_260_update_start_
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_260_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_260_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_273_update_start_
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_273_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_273_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_285_update_start_
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_285_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_285_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_298_update_start_
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_298_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_310_update_start_
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_310_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_310_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_323_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_335_update_start_
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_335_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_335_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_348_update_start_
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_348_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_348_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_360_update_start_
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_360_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_360_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_373_update_start_
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_373_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_373_Update/cr
      -- 
    rr_137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => RPIPE_ConvTranspose_input_pipe_28_inst_req_0); -- 
    cr_156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_32_inst_req_1); -- 
    cr_380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_132_inst_req_1); -- 
    cr_184_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_184_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_45_inst_req_1); -- 
    cr_212_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_212_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_57_inst_req_1); -- 
    cr_240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_70_inst_req_1); -- 
    cr_268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_82_inst_req_1); -- 
    cr_296_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_296_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_95_inst_req_1); -- 
    cr_324_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_324_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_107_inst_req_1); -- 
    cr_352_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_352_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_120_inst_req_1); -- 
    cr_408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_145_inst_req_1); -- 
    cr_436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_157_inst_req_1); -- 
    cr_464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_170_inst_req_1); -- 
    cr_492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_182_inst_req_1); -- 
    cr_520_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_520_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_195_inst_req_1); -- 
    cr_534_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_534_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_204_inst_req_1); -- 
    cr_548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_208_inst_req_1); -- 
    cr_562_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_562_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_212_inst_req_1); -- 
    cr_576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_226_inst_req_1); -- 
    cr_590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_230_inst_req_1); -- 
    cr_604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_234_inst_req_1); -- 
    cr_618_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_618_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_238_inst_req_1); -- 
    cr_646_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_646_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_260_inst_req_1); -- 
    cr_674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_273_inst_req_1); -- 
    cr_702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_285_inst_req_1); -- 
    cr_730_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_730_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_298_inst_req_1); -- 
    cr_758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_310_inst_req_1); -- 
    cr_786_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_786_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_323_inst_req_1); -- 
    cr_814_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_814_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_335_inst_req_1); -- 
    cr_842_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_842_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_348_inst_req_1); -- 
    cr_870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_360_inst_req_1); -- 
    cr_898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_373_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_28_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_28_update_start_
      -- CP-element group 1: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_28_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_28_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_28_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_28_Update/cr
      -- 
    ra_138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_28_inst_ack_0, ack => convTranspose_CP_39_elements(1)); -- 
    cr_142_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_142_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(1), ack => RPIPE_ConvTranspose_input_pipe_28_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_28_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_28_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_28_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_32_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_32_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_32_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_41_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_41_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_41_Sample/rr
      -- 
    ca_143_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_28_inst_ack_1, ack => convTranspose_CP_39_elements(2)); -- 
    rr_151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(2), ack => type_cast_32_inst_req_0); -- 
    rr_165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(2), ack => RPIPE_ConvTranspose_input_pipe_41_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_32_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_32_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_32_Sample/ra
      -- 
    ra_152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_32_inst_ack_0, ack => convTranspose_CP_39_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	57 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_32_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_32_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_32_Update/ca
      -- 
    ca_157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_32_inst_ack_1, ack => convTranspose_CP_39_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_41_Update/cr
      -- CP-element group 5: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_41_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_41_update_start_
      -- CP-element group 5: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_41_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_41_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_41_Update/$entry
      -- 
    ra_166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_41_inst_ack_0, ack => convTranspose_CP_39_elements(5)); -- 
    cr_170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(5), ack => RPIPE_ConvTranspose_input_pipe_41_inst_req_1); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_41_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_45_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_41_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_41_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_45_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_45_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_53_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_53_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_53_Sample/rr
      -- 
    ca_171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_41_inst_ack_1, ack => convTranspose_CP_39_elements(6)); -- 
    rr_179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(6), ack => type_cast_45_inst_req_0); -- 
    rr_193_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_193_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(6), ack => RPIPE_ConvTranspose_input_pipe_53_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_45_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_45_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_45_Sample/ra
      -- 
    ra_180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_45_inst_ack_0, ack => convTranspose_CP_39_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	57 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_45_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_45_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_45_Update/ca
      -- 
    ca_185_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_45_inst_ack_1, ack => convTranspose_CP_39_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_53_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_53_update_start_
      -- CP-element group 9: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_53_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_53_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_53_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_53_Update/cr
      -- 
    ra_194_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_53_inst_ack_0, ack => convTranspose_CP_39_elements(9)); -- 
    cr_198_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_198_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(9), ack => RPIPE_ConvTranspose_input_pipe_53_inst_req_1); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	13 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_53_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_53_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_53_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_57_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_57_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_57_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_66_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_66_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_66_Sample/rr
      -- 
    ca_199_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_53_inst_ack_1, ack => convTranspose_CP_39_elements(10)); -- 
    rr_207_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_207_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(10), ack => type_cast_57_inst_req_0); -- 
    rr_221_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_221_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(10), ack => RPIPE_ConvTranspose_input_pipe_66_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_57_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_57_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_57_Sample/ra
      -- 
    ra_208_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_57_inst_ack_0, ack => convTranspose_CP_39_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	60 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_57_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_57_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_57_Update/ca
      -- 
    ca_213_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_57_inst_ack_1, ack => convTranspose_CP_39_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_66_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_66_update_start_
      -- CP-element group 13: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_66_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_66_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_66_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_66_Update/cr
      -- 
    ra_222_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_66_inst_ack_0, ack => convTranspose_CP_39_elements(13)); -- 
    cr_226_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_226_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(13), ack => RPIPE_ConvTranspose_input_pipe_66_inst_req_1); -- 
    -- CP-element group 14:  fork  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_66_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_66_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_66_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_70_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_70_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_70_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_78_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_78_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_78_Sample/rr
      -- 
    ca_227_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_66_inst_ack_1, ack => convTranspose_CP_39_elements(14)); -- 
    rr_235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(14), ack => type_cast_70_inst_req_0); -- 
    rr_249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(14), ack => RPIPE_ConvTranspose_input_pipe_78_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_70_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_70_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_70_Sample/ra
      -- 
    ra_236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_70_inst_ack_0, ack => convTranspose_CP_39_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	0 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	60 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_70_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_70_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_70_Update/ca
      -- 
    ca_241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_70_inst_ack_1, ack => convTranspose_CP_39_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_78_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_78_update_start_
      -- CP-element group 17: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_78_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_78_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_78_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_78_Update/cr
      -- 
    ra_250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_78_inst_ack_0, ack => convTranspose_CP_39_elements(17)); -- 
    cr_254_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_254_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(17), ack => RPIPE_ConvTranspose_input_pipe_78_inst_req_1); -- 
    -- CP-element group 18:  fork  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18: 	21 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_78_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_78_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_78_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_82_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_82_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_82_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_91_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_91_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_91_Sample/rr
      -- 
    ca_255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_78_inst_ack_1, ack => convTranspose_CP_39_elements(18)); -- 
    rr_263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(18), ack => type_cast_82_inst_req_0); -- 
    rr_277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(18), ack => RPIPE_ConvTranspose_input_pipe_91_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_82_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_82_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_82_Sample/ra
      -- 
    ra_264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_82_inst_ack_0, ack => convTranspose_CP_39_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	63 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_82_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_82_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_82_Update/ca
      -- 
    ca_269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_82_inst_ack_1, ack => convTranspose_CP_39_elements(20)); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_91_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_91_update_start_
      -- CP-element group 21: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_91_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_91_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_91_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_91_Update/cr
      -- 
    ra_278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_91_inst_ack_0, ack => convTranspose_CP_39_elements(21)); -- 
    cr_282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(21), ack => RPIPE_ConvTranspose_input_pipe_91_inst_req_1); -- 
    -- CP-element group 22:  fork  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22: 	25 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_91_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_91_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_91_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_95_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_95_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_95_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_103_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_103_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_103_Sample/rr
      -- 
    ca_283_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_91_inst_ack_1, ack => convTranspose_CP_39_elements(22)); -- 
    rr_291_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_291_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(22), ack => type_cast_95_inst_req_0); -- 
    rr_305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(22), ack => RPIPE_ConvTranspose_input_pipe_103_inst_req_0); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_95_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_95_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_95_Sample/ra
      -- 
    ra_292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_95_inst_ack_0, ack => convTranspose_CP_39_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	0 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	63 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_95_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_95_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_95_Update/ca
      -- 
    ca_297_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_95_inst_ack_1, ack => convTranspose_CP_39_elements(24)); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	22 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_103_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_103_update_start_
      -- CP-element group 25: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_103_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_103_Sample/ra
      -- CP-element group 25: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_103_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_103_Update/cr
      -- 
    ra_306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_103_inst_ack_0, ack => convTranspose_CP_39_elements(25)); -- 
    cr_310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(25), ack => RPIPE_ConvTranspose_input_pipe_103_inst_req_1); -- 
    -- CP-element group 26:  fork  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: 	29 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_103_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_103_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_103_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_107_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_107_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_107_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_116_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_116_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_116_Sample/rr
      -- 
    ca_311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_103_inst_ack_1, ack => convTranspose_CP_39_elements(26)); -- 
    rr_319_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_319_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(26), ack => type_cast_107_inst_req_0); -- 
    rr_333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(26), ack => RPIPE_ConvTranspose_input_pipe_116_inst_req_0); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_107_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_107_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_107_Sample/ra
      -- 
    ra_320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_107_inst_ack_0, ack => convTranspose_CP_39_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	0 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	66 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_107_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_107_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_107_Update/ca
      -- 
    ca_325_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_107_inst_ack_1, ack => convTranspose_CP_39_elements(28)); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	26 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_116_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_116_update_start_
      -- CP-element group 29: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_116_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_116_Sample/ra
      -- CP-element group 29: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_116_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_116_Update/cr
      -- 
    ra_334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_116_inst_ack_0, ack => convTranspose_CP_39_elements(29)); -- 
    cr_338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(29), ack => RPIPE_ConvTranspose_input_pipe_116_inst_req_1); -- 
    -- CP-element group 30:  fork  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: 	33 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_116_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_116_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_116_Update/ca
      -- CP-element group 30: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_120_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_120_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_120_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_128_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_128_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_128_Sample/rr
      -- 
    ca_339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_116_inst_ack_1, ack => convTranspose_CP_39_elements(30)); -- 
    rr_347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(30), ack => type_cast_120_inst_req_0); -- 
    rr_361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(30), ack => RPIPE_ConvTranspose_input_pipe_128_inst_req_0); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_120_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_120_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_120_Sample/ra
      -- 
    ra_348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_120_inst_ack_0, ack => convTranspose_CP_39_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	0 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	66 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_120_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_120_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_120_Update/ca
      -- 
    ca_353_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_120_inst_ack_1, ack => convTranspose_CP_39_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	30 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_128_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_128_update_start_
      -- CP-element group 33: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_128_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_128_Sample/ra
      -- CP-element group 33: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_128_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_128_Update/cr
      -- 
    ra_362_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_128_inst_ack_0, ack => convTranspose_CP_39_elements(33)); -- 
    cr_366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(33), ack => RPIPE_ConvTranspose_input_pipe_128_inst_req_1); -- 
    -- CP-element group 34:  fork  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	37 
    -- CP-element group 34:  members (9) 
      -- CP-element group 34: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_132_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_132_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_132_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_128_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_128_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_128_Update/ca
      -- CP-element group 34: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_141_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_141_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_141_Sample/rr
      -- 
    ca_367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_128_inst_ack_1, ack => convTranspose_CP_39_elements(34)); -- 
    rr_375_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_375_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(34), ack => type_cast_132_inst_req_0); -- 
    rr_389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(34), ack => RPIPE_ConvTranspose_input_pipe_141_inst_req_0); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_132_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_132_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_132_Sample/ra
      -- 
    ra_376_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_132_inst_ack_0, ack => convTranspose_CP_39_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	0 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	69 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_132_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_132_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_132_Update/ca
      -- 
    ca_381_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_132_inst_ack_1, ack => convTranspose_CP_39_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_141_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_141_update_start_
      -- CP-element group 37: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_141_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_141_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_141_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_141_Update/cr
      -- 
    ra_390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_141_inst_ack_0, ack => convTranspose_CP_39_elements(37)); -- 
    cr_394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(37), ack => RPIPE_ConvTranspose_input_pipe_141_inst_req_1); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	41 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_141_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_141_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_141_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_145_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_145_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_145_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_153_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_153_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_153_Sample/rr
      -- 
    ca_395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_141_inst_ack_1, ack => convTranspose_CP_39_elements(38)); -- 
    rr_403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(38), ack => type_cast_145_inst_req_0); -- 
    rr_417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(38), ack => RPIPE_ConvTranspose_input_pipe_153_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_145_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_145_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_145_Sample/ra
      -- 
    ra_404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_145_inst_ack_0, ack => convTranspose_CP_39_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	0 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	69 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_145_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_145_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_145_Update/ca
      -- 
    ca_409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_145_inst_ack_1, ack => convTranspose_CP_39_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	38 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_153_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_153_update_start_
      -- CP-element group 41: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_153_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_153_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_153_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_153_Update/cr
      -- 
    ra_418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_153_inst_ack_0, ack => convTranspose_CP_39_elements(41)); -- 
    cr_422_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_422_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(41), ack => RPIPE_ConvTranspose_input_pipe_153_inst_req_1); -- 
    -- CP-element group 42:  fork  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	45 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (9) 
      -- CP-element group 42: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_153_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_153_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_153_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_157_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_157_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_157_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_166_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_166_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_166_Sample/rr
      -- 
    ca_423_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_153_inst_ack_1, ack => convTranspose_CP_39_elements(42)); -- 
    rr_445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(42), ack => RPIPE_ConvTranspose_input_pipe_166_inst_req_0); -- 
    rr_431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(42), ack => type_cast_157_inst_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_157_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_157_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_157_Sample/ra
      -- 
    ra_432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_157_inst_ack_0, ack => convTranspose_CP_39_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	0 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	72 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_157_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_157_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_157_Update/ca
      -- 
    ca_437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_157_inst_ack_1, ack => convTranspose_CP_39_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	42 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_166_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_166_update_start_
      -- CP-element group 45: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_166_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_166_Sample/ra
      -- CP-element group 45: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_166_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_166_Update/cr
      -- 
    ra_446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_166_inst_ack_0, ack => convTranspose_CP_39_elements(45)); -- 
    cr_450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(45), ack => RPIPE_ConvTranspose_input_pipe_166_inst_req_1); -- 
    -- CP-element group 46:  fork  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46: 	49 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_166_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_166_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_166_Update/ca
      -- CP-element group 46: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_170_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_170_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_170_Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_178_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_178_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_178_Sample/rr
      -- 
    ca_451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_166_inst_ack_1, ack => convTranspose_CP_39_elements(46)); -- 
    rr_459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(46), ack => type_cast_170_inst_req_0); -- 
    rr_473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(46), ack => RPIPE_ConvTranspose_input_pipe_178_inst_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_170_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_170_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_170_Sample/ra
      -- 
    ra_460_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_170_inst_ack_0, ack => convTranspose_CP_39_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	0 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	72 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_170_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_170_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_170_Update/ca
      -- 
    ca_465_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_170_inst_ack_1, ack => convTranspose_CP_39_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	46 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_178_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_178_update_start_
      -- CP-element group 49: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_178_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_178_Sample/ra
      -- CP-element group 49: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_178_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_178_Update/cr
      -- 
    ra_474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_178_inst_ack_0, ack => convTranspose_CP_39_elements(49)); -- 
    cr_478_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_478_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(49), ack => RPIPE_ConvTranspose_input_pipe_178_inst_req_1); -- 
    -- CP-element group 50:  fork  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	53 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_178_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_178_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_178_Update/ca
      -- CP-element group 50: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_182_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_182_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_182_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_191_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_191_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_191_Sample/rr
      -- 
    ca_479_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_178_inst_ack_1, ack => convTranspose_CP_39_elements(50)); -- 
    rr_487_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_487_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(50), ack => type_cast_182_inst_req_0); -- 
    rr_501_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_501_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(50), ack => RPIPE_ConvTranspose_input_pipe_191_inst_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_182_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_182_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_182_Sample/ra
      -- 
    ra_488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_182_inst_ack_0, ack => convTranspose_CP_39_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	0 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	75 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_182_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_182_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_182_Update/ca
      -- 
    ca_493_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_182_inst_ack_1, ack => convTranspose_CP_39_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	50 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (6) 
      -- CP-element group 53: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_191_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_191_update_start_
      -- CP-element group 53: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_191_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_191_Sample/ra
      -- CP-element group 53: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_191_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_191_Update/cr
      -- 
    ra_502_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_191_inst_ack_0, ack => convTranspose_CP_39_elements(53)); -- 
    cr_506_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_506_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(53), ack => RPIPE_ConvTranspose_input_pipe_191_inst_req_1); -- 
    -- CP-element group 54:  fork  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54: 	78 
    -- CP-element group 54:  members (9) 
      -- CP-element group 54: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_191_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_191_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_191_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_195_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_195_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_195_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_256_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_256_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_256_Sample/rr
      -- 
    ca_507_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_191_inst_ack_1, ack => convTranspose_CP_39_elements(54)); -- 
    rr_515_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_515_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(54), ack => type_cast_195_inst_req_0); -- 
    rr_627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(54), ack => RPIPE_ConvTranspose_input_pipe_256_inst_req_0); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_195_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_195_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_195_Sample/ra
      -- 
    ra_516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_195_inst_ack_0, ack => convTranspose_CP_39_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	0 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	75 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_195_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_195_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_195_Update/ca
      -- 
    ca_521_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_195_inst_ack_1, ack => convTranspose_CP_39_elements(56)); -- 
    -- CP-element group 57:  join  transition  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	4 
    -- CP-element group 57: 	8 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_204_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_204_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_204_Sample/rr
      -- 
    rr_529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(57), ack => type_cast_204_inst_req_0); -- 
    convTranspose_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(4) & convTranspose_CP_39_elements(8);
      gj_convTranspose_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_204_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_204_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_204_Sample/ra
      -- 
    ra_530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_204_inst_ack_0, ack => convTranspose_CP_39_elements(58)); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	0 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	118 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_204_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_204_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_204_Update/ca
      -- 
    ca_535_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_204_inst_ack_1, ack => convTranspose_CP_39_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	12 
    -- CP-element group 60: 	16 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_208_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_208_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_208_Sample/rr
      -- 
    rr_543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(60), ack => type_cast_208_inst_req_0); -- 
    convTranspose_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(12) & convTranspose_CP_39_elements(16);
      gj_convTranspose_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_208_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_208_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_208_Sample/ra
      -- 
    ra_544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_208_inst_ack_0, ack => convTranspose_CP_39_elements(61)); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	0 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	118 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_208_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_208_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_208_Update/ca
      -- 
    ca_549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_208_inst_ack_1, ack => convTranspose_CP_39_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	20 
    -- CP-element group 63: 	24 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_212_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_212_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_212_Sample/rr
      -- 
    rr_557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(63), ack => type_cast_212_inst_req_0); -- 
    convTranspose_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(20) & convTranspose_CP_39_elements(24);
      gj_convTranspose_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_212_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_212_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_212_Sample/ra
      -- 
    ra_558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_212_inst_ack_0, ack => convTranspose_CP_39_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	0 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	118 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_212_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_212_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_212_Update/ca
      -- 
    ca_563_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_212_inst_ack_1, ack => convTranspose_CP_39_elements(65)); -- 
    -- CP-element group 66:  join  transition  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	28 
    -- CP-element group 66: 	32 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_226_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_226_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_226_Sample/rr
      -- 
    rr_571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(66), ack => type_cast_226_inst_req_0); -- 
    convTranspose_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(28) & convTranspose_CP_39_elements(32);
      gj_convTranspose_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_226_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_226_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_226_Sample/ra
      -- 
    ra_572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_226_inst_ack_0, ack => convTranspose_CP_39_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	0 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	118 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_226_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_226_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_226_Update/ca
      -- 
    ca_577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_226_inst_ack_1, ack => convTranspose_CP_39_elements(68)); -- 
    -- CP-element group 69:  join  transition  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	40 
    -- CP-element group 69: 	36 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_230_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_230_Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_230_Sample/rr
      -- 
    rr_585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(69), ack => type_cast_230_inst_req_0); -- 
    convTranspose_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(40) & convTranspose_CP_39_elements(36);
      gj_convTranspose_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_230_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_230_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_230_Sample/ra
      -- 
    ra_586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_230_inst_ack_0, ack => convTranspose_CP_39_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	0 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	118 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_230_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_230_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_230_Update/ca
      -- 
    ca_591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_230_inst_ack_1, ack => convTranspose_CP_39_elements(71)); -- 
    -- CP-element group 72:  join  transition  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	44 
    -- CP-element group 72: 	48 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_234_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_234_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_234_Sample/rr
      -- 
    rr_599_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_599_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(72), ack => type_cast_234_inst_req_0); -- 
    convTranspose_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(44) & convTranspose_CP_39_elements(48);
      gj_convTranspose_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_234_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_234_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_234_Sample/ra
      -- 
    ra_600_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_234_inst_ack_0, ack => convTranspose_CP_39_elements(73)); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	0 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	118 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_234_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_234_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_234_Update/ca
      -- 
    ca_605_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_234_inst_ack_1, ack => convTranspose_CP_39_elements(74)); -- 
    -- CP-element group 75:  join  transition  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	56 
    -- CP-element group 75: 	52 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_238_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_238_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_238_Sample/rr
      -- 
    rr_613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(75), ack => type_cast_238_inst_req_0); -- 
    convTranspose_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(56) & convTranspose_CP_39_elements(52);
      gj_convTranspose_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_238_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_238_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_238_Sample/ra
      -- 
    ra_614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_238_inst_ack_0, ack => convTranspose_CP_39_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	0 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	118 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_238_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_238_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_238_Update/ca
      -- 
    ca_619_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_238_inst_ack_1, ack => convTranspose_CP_39_elements(77)); -- 
    -- CP-element group 78:  transition  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	54 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (6) 
      -- CP-element group 78: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_256_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_256_update_start_
      -- CP-element group 78: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_256_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_256_Sample/ra
      -- CP-element group 78: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_256_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_256_Update/cr
      -- 
    ra_628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_256_inst_ack_0, ack => convTranspose_CP_39_elements(78)); -- 
    cr_632_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_632_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(78), ack => RPIPE_ConvTranspose_input_pipe_256_inst_req_1); -- 
    -- CP-element group 79:  fork  transition  input  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79: 	82 
    -- CP-element group 79:  members (9) 
      -- CP-element group 79: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_256_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_256_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_256_Update/ca
      -- CP-element group 79: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_260_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_260_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_260_Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_269_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_269_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_269_Sample/rr
      -- 
    ca_633_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_256_inst_ack_1, ack => convTranspose_CP_39_elements(79)); -- 
    rr_641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(79), ack => type_cast_260_inst_req_0); -- 
    rr_655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(79), ack => RPIPE_ConvTranspose_input_pipe_269_inst_req_0); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_260_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_260_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_260_Sample/ra
      -- 
    ra_642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_260_inst_ack_0, ack => convTranspose_CP_39_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	0 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	118 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_260_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_260_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_260_Update/ca
      -- 
    ca_647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_260_inst_ack_1, ack => convTranspose_CP_39_elements(81)); -- 
    -- CP-element group 82:  transition  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	79 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (6) 
      -- CP-element group 82: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_269_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_269_update_start_
      -- CP-element group 82: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_269_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_269_Sample/ra
      -- CP-element group 82: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_269_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_269_Update/cr
      -- 
    ra_656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_269_inst_ack_0, ack => convTranspose_CP_39_elements(82)); -- 
    cr_660_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_660_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(82), ack => RPIPE_ConvTranspose_input_pipe_269_inst_req_1); -- 
    -- CP-element group 83:  fork  transition  input  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83: 	86 
    -- CP-element group 83:  members (9) 
      -- CP-element group 83: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_269_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_269_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_269_Update/ca
      -- CP-element group 83: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_273_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_273_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_273_Sample/rr
      -- CP-element group 83: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_281_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_281_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_281_Sample/rr
      -- 
    ca_661_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_269_inst_ack_1, ack => convTranspose_CP_39_elements(83)); -- 
    rr_669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(83), ack => type_cast_273_inst_req_0); -- 
    rr_683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(83), ack => RPIPE_ConvTranspose_input_pipe_281_inst_req_0); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_273_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_273_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_273_Sample/ra
      -- 
    ra_670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_273_inst_ack_0, ack => convTranspose_CP_39_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	0 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	118 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_273_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_273_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_273_Update/ca
      -- 
    ca_675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_273_inst_ack_1, ack => convTranspose_CP_39_elements(85)); -- 
    -- CP-element group 86:  transition  input  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	83 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (6) 
      -- CP-element group 86: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_281_sample_completed_
      -- CP-element group 86: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_281_update_start_
      -- CP-element group 86: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_281_Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_281_Sample/ra
      -- CP-element group 86: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_281_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_281_Update/cr
      -- 
    ra_684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_281_inst_ack_0, ack => convTranspose_CP_39_elements(86)); -- 
    cr_688_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_688_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(86), ack => RPIPE_ConvTranspose_input_pipe_281_inst_req_1); -- 
    -- CP-element group 87:  fork  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87: 	90 
    -- CP-element group 87:  members (9) 
      -- CP-element group 87: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_281_update_completed_
      -- CP-element group 87: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_281_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_281_Update/ca
      -- CP-element group 87: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_285_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_285_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_285_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_294_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_294_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_294_Sample/rr
      -- 
    ca_689_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_281_inst_ack_1, ack => convTranspose_CP_39_elements(87)); -- 
    rr_697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(87), ack => type_cast_285_inst_req_0); -- 
    rr_711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(87), ack => RPIPE_ConvTranspose_input_pipe_294_inst_req_0); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_285_sample_completed_
      -- CP-element group 88: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_285_Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_285_Sample/ra
      -- 
    ra_698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_285_inst_ack_0, ack => convTranspose_CP_39_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	0 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	118 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_285_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_285_Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_285_Update/ca
      -- 
    ca_703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_285_inst_ack_1, ack => convTranspose_CP_39_elements(89)); -- 
    -- CP-element group 90:  transition  input  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	87 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (6) 
      -- CP-element group 90: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_294_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_294_update_start_
      -- CP-element group 90: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_294_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_294_Sample/ra
      -- CP-element group 90: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_294_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_294_Update/cr
      -- 
    ra_712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_294_inst_ack_0, ack => convTranspose_CP_39_elements(90)); -- 
    cr_716_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_716_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(90), ack => RPIPE_ConvTranspose_input_pipe_294_inst_req_1); -- 
    -- CP-element group 91:  fork  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91: 	94 
    -- CP-element group 91:  members (9) 
      -- CP-element group 91: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_294_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_294_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_294_Update/ca
      -- CP-element group 91: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_298_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_298_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_298_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_306_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_306_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_306_Sample/rr
      -- 
    ca_717_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_294_inst_ack_1, ack => convTranspose_CP_39_elements(91)); -- 
    rr_725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(91), ack => type_cast_298_inst_req_0); -- 
    rr_739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(91), ack => RPIPE_ConvTranspose_input_pipe_306_inst_req_0); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_298_sample_completed_
      -- CP-element group 92: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_298_Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_298_Sample/ra
      -- 
    ra_726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_298_inst_ack_0, ack => convTranspose_CP_39_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	0 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	118 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_298_Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_298_update_completed_
      -- CP-element group 93: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_298_Update/ca
      -- 
    ca_731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_298_inst_ack_1, ack => convTranspose_CP_39_elements(93)); -- 
    -- CP-element group 94:  transition  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	91 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (6) 
      -- CP-element group 94: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_306_sample_completed_
      -- CP-element group 94: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_306_update_start_
      -- CP-element group 94: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_306_Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_306_Sample/ra
      -- CP-element group 94: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_306_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_306_Update/cr
      -- 
    ra_740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_306_inst_ack_0, ack => convTranspose_CP_39_elements(94)); -- 
    cr_744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(94), ack => RPIPE_ConvTranspose_input_pipe_306_inst_req_1); -- 
    -- CP-element group 95:  fork  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95: 	98 
    -- CP-element group 95:  members (9) 
      -- CP-element group 95: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_319_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_319_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_319_Sample/rr
      -- CP-element group 95: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_306_update_completed_
      -- CP-element group 95: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_306_Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_306_Update/ca
      -- CP-element group 95: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_310_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_310_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_310_Sample/rr
      -- 
    ca_745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_306_inst_ack_1, ack => convTranspose_CP_39_elements(95)); -- 
    rr_753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(95), ack => type_cast_310_inst_req_0); -- 
    rr_767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(95), ack => RPIPE_ConvTranspose_input_pipe_319_inst_req_0); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_310_sample_completed_
      -- CP-element group 96: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_310_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_310_Sample/ra
      -- 
    ra_754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_310_inst_ack_0, ack => convTranspose_CP_39_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	0 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	118 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_310_update_completed_
      -- CP-element group 97: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_310_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_310_Update/ca
      -- 
    ca_759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_310_inst_ack_1, ack => convTranspose_CP_39_elements(97)); -- 
    -- CP-element group 98:  transition  input  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	95 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (6) 
      -- CP-element group 98: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_319_sample_completed_
      -- CP-element group 98: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_319_update_start_
      -- CP-element group 98: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_319_Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_319_Sample/ra
      -- CP-element group 98: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_319_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_319_Update/cr
      -- 
    ra_768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_319_inst_ack_0, ack => convTranspose_CP_39_elements(98)); -- 
    cr_772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(98), ack => RPIPE_ConvTranspose_input_pipe_319_inst_req_1); -- 
    -- CP-element group 99:  fork  transition  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: 	102 
    -- CP-element group 99:  members (9) 
      -- CP-element group 99: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_319_update_completed_
      -- CP-element group 99: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_319_Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_319_Update/ca
      -- CP-element group 99: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_323_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_323_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_323_Sample/rr
      -- CP-element group 99: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_331_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_331_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_331_Sample/rr
      -- 
    ca_773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_319_inst_ack_1, ack => convTranspose_CP_39_elements(99)); -- 
    rr_781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(99), ack => type_cast_323_inst_req_0); -- 
    rr_795_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_795_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(99), ack => RPIPE_ConvTranspose_input_pipe_331_inst_req_0); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_323_sample_completed_
      -- CP-element group 100: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_323_Sample/$exit
      -- CP-element group 100: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_323_Sample/ra
      -- 
    ra_782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_323_inst_ack_0, ack => convTranspose_CP_39_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	0 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	118 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_323_update_completed_
      -- CP-element group 101: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_323_Update/$exit
      -- CP-element group 101: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_323_Update/ca
      -- 
    ca_787_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_323_inst_ack_1, ack => convTranspose_CP_39_elements(101)); -- 
    -- CP-element group 102:  transition  input  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	99 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102:  members (6) 
      -- CP-element group 102: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_331_sample_completed_
      -- CP-element group 102: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_331_update_start_
      -- CP-element group 102: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_331_Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_331_Sample/ra
      -- CP-element group 102: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_331_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_331_Update/cr
      -- 
    ra_796_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_331_inst_ack_0, ack => convTranspose_CP_39_elements(102)); -- 
    cr_800_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_800_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(102), ack => RPIPE_ConvTranspose_input_pipe_331_inst_req_1); -- 
    -- CP-element group 103:  fork  transition  input  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103: 	106 
    -- CP-element group 103:  members (9) 
      -- CP-element group 103: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_331_update_completed_
      -- CP-element group 103: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_331_Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_331_Update/ca
      -- CP-element group 103: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_335_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_335_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_335_Sample/rr
      -- CP-element group 103: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_344_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_344_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_344_Sample/rr
      -- 
    ca_801_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_331_inst_ack_1, ack => convTranspose_CP_39_elements(103)); -- 
    rr_809_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_809_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(103), ack => type_cast_335_inst_req_0); -- 
    rr_823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(103), ack => RPIPE_ConvTranspose_input_pipe_344_inst_req_0); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_335_sample_completed_
      -- CP-element group 104: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_335_Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_335_Sample/ra
      -- 
    ra_810_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_335_inst_ack_0, ack => convTranspose_CP_39_elements(104)); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	0 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	118 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_335_update_completed_
      -- CP-element group 105: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_335_Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_335_Update/ca
      -- 
    ca_815_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_335_inst_ack_1, ack => convTranspose_CP_39_elements(105)); -- 
    -- CP-element group 106:  transition  input  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	103 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (6) 
      -- CP-element group 106: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_344_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_344_update_start_
      -- CP-element group 106: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_344_Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_344_Sample/ra
      -- CP-element group 106: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_344_Update/$entry
      -- CP-element group 106: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_344_Update/cr
      -- 
    ra_824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_344_inst_ack_0, ack => convTranspose_CP_39_elements(106)); -- 
    cr_828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(106), ack => RPIPE_ConvTranspose_input_pipe_344_inst_req_1); -- 
    -- CP-element group 107:  fork  transition  input  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107: 	110 
    -- CP-element group 107:  members (9) 
      -- CP-element group 107: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_344_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_344_Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_344_Update/ca
      -- CP-element group 107: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_348_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_348_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_348_Sample/rr
      -- CP-element group 107: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_356_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_356_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_356_Sample/rr
      -- 
    ca_829_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_344_inst_ack_1, ack => convTranspose_CP_39_elements(107)); -- 
    rr_837_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_837_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(107), ack => type_cast_348_inst_req_0); -- 
    rr_851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(107), ack => RPIPE_ConvTranspose_input_pipe_356_inst_req_0); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_348_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_348_Sample/$exit
      -- CP-element group 108: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_348_Sample/ra
      -- 
    ra_838_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_348_inst_ack_0, ack => convTranspose_CP_39_elements(108)); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	0 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	118 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_348_update_completed_
      -- CP-element group 109: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_348_Update/$exit
      -- CP-element group 109: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_348_Update/ca
      -- 
    ca_843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_348_inst_ack_1, ack => convTranspose_CP_39_elements(109)); -- 
    -- CP-element group 110:  transition  input  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	107 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (6) 
      -- CP-element group 110: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_356_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_356_update_start_
      -- CP-element group 110: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_356_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_356_Sample/ra
      -- CP-element group 110: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_356_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_356_Update/cr
      -- 
    ra_852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_356_inst_ack_0, ack => convTranspose_CP_39_elements(110)); -- 
    cr_856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(110), ack => RPIPE_ConvTranspose_input_pipe_356_inst_req_1); -- 
    -- CP-element group 111:  fork  transition  input  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111: 	114 
    -- CP-element group 111:  members (9) 
      -- CP-element group 111: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_356_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_356_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_356_Update/ca
      -- CP-element group 111: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_360_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_360_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_360_Sample/rr
      -- CP-element group 111: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_369_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_369_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_369_Sample/rr
      -- 
    ca_857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_356_inst_ack_1, ack => convTranspose_CP_39_elements(111)); -- 
    rr_865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(111), ack => type_cast_360_inst_req_0); -- 
    rr_879_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_879_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(111), ack => RPIPE_ConvTranspose_input_pipe_369_inst_req_0); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_360_sample_completed_
      -- CP-element group 112: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_360_Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_360_Sample/ra
      -- 
    ra_866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_360_inst_ack_0, ack => convTranspose_CP_39_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	0 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	118 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_360_update_completed_
      -- CP-element group 113: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_360_Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_360_Update/ca
      -- 
    ca_871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_360_inst_ack_1, ack => convTranspose_CP_39_elements(113)); -- 
    -- CP-element group 114:  transition  input  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	111 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (6) 
      -- CP-element group 114: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_369_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_369_update_start_
      -- CP-element group 114: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_369_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_369_Sample/ra
      -- CP-element group 114: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_369_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_369_Update/cr
      -- 
    ra_880_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_369_inst_ack_0, ack => convTranspose_CP_39_elements(114)); -- 
    cr_884_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_884_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(114), ack => RPIPE_ConvTranspose_input_pipe_369_inst_req_1); -- 
    -- CP-element group 115:  transition  input  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (6) 
      -- CP-element group 115: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_369_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_369_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/RPIPE_ConvTranspose_input_pipe_369_Update/ca
      -- CP-element group 115: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_373_sample_start_
      -- CP-element group 115: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_373_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_373_Sample/rr
      -- 
    ca_885_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_369_inst_ack_1, ack => convTranspose_CP_39_elements(115)); -- 
    rr_893_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_893_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(115), ack => type_cast_373_inst_req_0); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_373_sample_completed_
      -- CP-element group 116: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_373_Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_373_Sample/ra
      -- 
    ra_894_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_373_inst_ack_0, ack => convTranspose_CP_39_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	0 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_373_update_completed_
      -- CP-element group 117: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_373_Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/type_cast_373_Update/ca
      -- 
    ca_899_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_373_inst_ack_1, ack => convTranspose_CP_39_elements(117)); -- 
    -- CP-element group 118:  branch  join  transition  place  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	59 
    -- CP-element group 118: 	62 
    -- CP-element group 118: 	65 
    -- CP-element group 118: 	68 
    -- CP-element group 118: 	71 
    -- CP-element group 118: 	74 
    -- CP-element group 118: 	77 
    -- CP-element group 118: 	81 
    -- CP-element group 118: 	85 
    -- CP-element group 118: 	89 
    -- CP-element group 118: 	93 
    -- CP-element group 118: 	97 
    -- CP-element group 118: 	101 
    -- CP-element group 118: 	105 
    -- CP-element group 118: 	109 
    -- CP-element group 118: 	113 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118: 	120 
    -- CP-element group 118:  members (10) 
      -- CP-element group 118: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386__exit__
      -- CP-element group 118: 	 branch_block_stmt_26/if_stmt_387__entry__
      -- CP-element group 118: 	 branch_block_stmt_26/assign_stmt_29_to_assign_stmt_386/$exit
      -- CP-element group 118: 	 branch_block_stmt_26/if_stmt_387_dead_link/$entry
      -- CP-element group 118: 	 branch_block_stmt_26/if_stmt_387_eval_test/$entry
      -- CP-element group 118: 	 branch_block_stmt_26/if_stmt_387_eval_test/$exit
      -- CP-element group 118: 	 branch_block_stmt_26/if_stmt_387_eval_test/branch_req
      -- CP-element group 118: 	 branch_block_stmt_26/R_cmp456_388_place
      -- CP-element group 118: 	 branch_block_stmt_26/if_stmt_387_if_link/$entry
      -- CP-element group 118: 	 branch_block_stmt_26/if_stmt_387_else_link/$entry
      -- 
    branch_req_907_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_907_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(118), ack => if_stmt_387_branch_req_0); -- 
    convTranspose_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(59) & convTranspose_CP_39_elements(62) & convTranspose_CP_39_elements(65) & convTranspose_CP_39_elements(68) & convTranspose_CP_39_elements(71) & convTranspose_CP_39_elements(74) & convTranspose_CP_39_elements(77) & convTranspose_CP_39_elements(81) & convTranspose_CP_39_elements(85) & convTranspose_CP_39_elements(89) & convTranspose_CP_39_elements(93) & convTranspose_CP_39_elements(97) & convTranspose_CP_39_elements(101) & convTranspose_CP_39_elements(105) & convTranspose_CP_39_elements(109) & convTranspose_CP_39_elements(113) & convTranspose_CP_39_elements(117);
      gj_convTranspose_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	123 
    -- CP-element group 119: 	124 
    -- CP-element group 119:  members (18) 
      -- CP-element group 119: 	 branch_block_stmt_26/merge_stmt_408__exit__
      -- CP-element group 119: 	 branch_block_stmt_26/assign_stmt_414_to_assign_stmt_443__entry__
      -- CP-element group 119: 	 branch_block_stmt_26/if_stmt_387_if_link/$exit
      -- CP-element group 119: 	 branch_block_stmt_26/if_stmt_387_if_link/if_choice_transition
      -- CP-element group 119: 	 branch_block_stmt_26/entry_bbx_xnph458
      -- CP-element group 119: 	 branch_block_stmt_26/assign_stmt_414_to_assign_stmt_443/$entry
      -- CP-element group 119: 	 branch_block_stmt_26/assign_stmt_414_to_assign_stmt_443/type_cast_429_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_26/assign_stmt_414_to_assign_stmt_443/type_cast_429_update_start_
      -- CP-element group 119: 	 branch_block_stmt_26/assign_stmt_414_to_assign_stmt_443/type_cast_429_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_26/assign_stmt_414_to_assign_stmt_443/type_cast_429_Sample/rr
      -- CP-element group 119: 	 branch_block_stmt_26/assign_stmt_414_to_assign_stmt_443/type_cast_429_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_26/assign_stmt_414_to_assign_stmt_443/type_cast_429_Update/cr
      -- CP-element group 119: 	 branch_block_stmt_26/entry_bbx_xnph458_PhiReq/$entry
      -- CP-element group 119: 	 branch_block_stmt_26/entry_bbx_xnph458_PhiReq/$exit
      -- CP-element group 119: 	 branch_block_stmt_26/merge_stmt_408_PhiReqMerge
      -- CP-element group 119: 	 branch_block_stmt_26/merge_stmt_408_PhiAck/$entry
      -- CP-element group 119: 	 branch_block_stmt_26/merge_stmt_408_PhiAck/$exit
      -- CP-element group 119: 	 branch_block_stmt_26/merge_stmt_408_PhiAck/dummy
      -- 
    if_choice_transition_912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_387_branch_ack_1, ack => convTranspose_CP_39_elements(119)); -- 
    rr_951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(119), ack => type_cast_429_inst_req_0); -- 
    cr_956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(119), ack => type_cast_429_inst_req_1); -- 
    -- CP-element group 120:  transition  place  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	118 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	360 
    -- CP-element group 120:  members (5) 
      -- CP-element group 120: 	 branch_block_stmt_26/if_stmt_387_else_link/$exit
      -- CP-element group 120: 	 branch_block_stmt_26/if_stmt_387_else_link/else_choice_transition
      -- CP-element group 120: 	 branch_block_stmt_26/entry_forx_xcond190x_xpreheader
      -- CP-element group 120: 	 branch_block_stmt_26/entry_forx_xcond190x_xpreheader_PhiReq/$entry
      -- CP-element group 120: 	 branch_block_stmt_26/entry_forx_xcond190x_xpreheader_PhiReq/$exit
      -- 
    else_choice_transition_916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_387_branch_ack_0, ack => convTranspose_CP_39_elements(120)); -- 
    -- CP-element group 121:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	360 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	167 
    -- CP-element group 121: 	168 
    -- CP-element group 121:  members (18) 
      -- CP-element group 121: 	 branch_block_stmt_26/merge_stmt_615__exit__
      -- CP-element group 121: 	 branch_block_stmt_26/assign_stmt_621_to_assign_stmt_650__entry__
      -- CP-element group 121: 	 branch_block_stmt_26/assign_stmt_621_to_assign_stmt_650/type_cast_636_Update/cr
      -- CP-element group 121: 	 branch_block_stmt_26/assign_stmt_621_to_assign_stmt_650/type_cast_636_Update/$entry
      -- CP-element group 121: 	 branch_block_stmt_26/assign_stmt_621_to_assign_stmt_650/type_cast_636_Sample/rr
      -- CP-element group 121: 	 branch_block_stmt_26/assign_stmt_621_to_assign_stmt_650/type_cast_636_Sample/$entry
      -- CP-element group 121: 	 branch_block_stmt_26/assign_stmt_621_to_assign_stmt_650/type_cast_636_update_start_
      -- CP-element group 121: 	 branch_block_stmt_26/assign_stmt_621_to_assign_stmt_650/type_cast_636_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_26/assign_stmt_621_to_assign_stmt_650/$entry
      -- CP-element group 121: 	 branch_block_stmt_26/if_stmt_402_if_link/$exit
      -- CP-element group 121: 	 branch_block_stmt_26/if_stmt_402_if_link/if_choice_transition
      -- CP-element group 121: 	 branch_block_stmt_26/forx_xcond190x_xpreheader_bbx_xnph454
      -- CP-element group 121: 	 branch_block_stmt_26/forx_xcond190x_xpreheader_bbx_xnph454_PhiReq/$entry
      -- CP-element group 121: 	 branch_block_stmt_26/forx_xcond190x_xpreheader_bbx_xnph454_PhiReq/$exit
      -- CP-element group 121: 	 branch_block_stmt_26/merge_stmt_615_PhiReqMerge
      -- CP-element group 121: 	 branch_block_stmt_26/merge_stmt_615_PhiAck/$entry
      -- CP-element group 121: 	 branch_block_stmt_26/merge_stmt_615_PhiAck/$exit
      -- CP-element group 121: 	 branch_block_stmt_26/merge_stmt_615_PhiAck/dummy
      -- 
    if_choice_transition_934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_402_branch_ack_1, ack => convTranspose_CP_39_elements(121)); -- 
    cr_1315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(121), ack => type_cast_636_inst_req_1); -- 
    rr_1310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(121), ack => type_cast_636_inst_req_0); -- 
    -- CP-element group 122:  transition  place  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	360 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	373 
    -- CP-element group 122:  members (5) 
      -- CP-element group 122: 	 branch_block_stmt_26/if_stmt_402_else_link/$exit
      -- CP-element group 122: 	 branch_block_stmt_26/if_stmt_402_else_link/else_choice_transition
      -- CP-element group 122: 	 branch_block_stmt_26/forx_xcond190x_xpreheader_forx_xend250
      -- CP-element group 122: 	 branch_block_stmt_26/forx_xcond190x_xpreheader_forx_xend250_PhiReq/$entry
      -- CP-element group 122: 	 branch_block_stmt_26/forx_xcond190x_xpreheader_forx_xend250_PhiReq/$exit
      -- 
    else_choice_transition_938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_402_branch_ack_0, ack => convTranspose_CP_39_elements(122)); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	119 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_26/assign_stmt_414_to_assign_stmt_443/type_cast_429_sample_completed_
      -- CP-element group 123: 	 branch_block_stmt_26/assign_stmt_414_to_assign_stmt_443/type_cast_429_Sample/$exit
      -- CP-element group 123: 	 branch_block_stmt_26/assign_stmt_414_to_assign_stmt_443/type_cast_429_Sample/ra
      -- 
    ra_952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_429_inst_ack_0, ack => convTranspose_CP_39_elements(123)); -- 
    -- CP-element group 124:  transition  place  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	119 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	361 
    -- CP-element group 124:  members (9) 
      -- CP-element group 124: 	 branch_block_stmt_26/assign_stmt_414_to_assign_stmt_443__exit__
      -- CP-element group 124: 	 branch_block_stmt_26/bbx_xnph458_forx_xbody
      -- CP-element group 124: 	 branch_block_stmt_26/assign_stmt_414_to_assign_stmt_443/$exit
      -- CP-element group 124: 	 branch_block_stmt_26/assign_stmt_414_to_assign_stmt_443/type_cast_429_update_completed_
      -- CP-element group 124: 	 branch_block_stmt_26/assign_stmt_414_to_assign_stmt_443/type_cast_429_Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_26/assign_stmt_414_to_assign_stmt_443/type_cast_429_Update/ca
      -- CP-element group 124: 	 branch_block_stmt_26/bbx_xnph458_forx_xbody_PhiReq/$entry
      -- CP-element group 124: 	 branch_block_stmt_26/bbx_xnph458_forx_xbody_PhiReq/phi_stmt_446/$entry
      -- CP-element group 124: 	 branch_block_stmt_26/bbx_xnph458_forx_xbody_PhiReq/phi_stmt_446/phi_stmt_446_sources/$entry
      -- 
    ca_957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_429_inst_ack_1, ack => convTranspose_CP_39_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	366 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	164 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/array_obj_ref_458_final_index_sum_regn_sample_complete
      -- CP-element group 125: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/array_obj_ref_458_final_index_sum_regn_Sample/$exit
      -- CP-element group 125: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/array_obj_ref_458_final_index_sum_regn_Sample/ack
      -- 
    ack_986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_458_index_offset_ack_0, ack => convTranspose_CP_39_elements(125)); -- 
    -- CP-element group 126:  transition  input  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	366 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (11) 
      -- CP-element group 126: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/addr_of_459_sample_start_
      -- CP-element group 126: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/array_obj_ref_458_root_address_calculated
      -- CP-element group 126: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/array_obj_ref_458_offset_calculated
      -- CP-element group 126: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/array_obj_ref_458_final_index_sum_regn_Update/$exit
      -- CP-element group 126: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/array_obj_ref_458_final_index_sum_regn_Update/ack
      -- CP-element group 126: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/array_obj_ref_458_base_plus_offset/$entry
      -- CP-element group 126: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/array_obj_ref_458_base_plus_offset/$exit
      -- CP-element group 126: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/array_obj_ref_458_base_plus_offset/sum_rename_req
      -- CP-element group 126: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/array_obj_ref_458_base_plus_offset/sum_rename_ack
      -- CP-element group 126: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/addr_of_459_request/$entry
      -- CP-element group 126: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/addr_of_459_request/req
      -- 
    ack_991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_458_index_offset_ack_1, ack => convTranspose_CP_39_elements(126)); -- 
    req_1000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(126), ack => addr_of_459_final_reg_req_0); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/addr_of_459_sample_completed_
      -- CP-element group 127: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/addr_of_459_request/$exit
      -- CP-element group 127: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/addr_of_459_request/ack
      -- 
    ack_1001_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_459_final_reg_ack_0, ack => convTranspose_CP_39_elements(127)); -- 
    -- CP-element group 128:  fork  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	366 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	161 
    -- CP-element group 128:  members (19) 
      -- CP-element group 128: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/ptr_deref_595_root_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/ptr_deref_595_base_address_resized
      -- CP-element group 128: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/ptr_deref_595_word_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/ptr_deref_595_base_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/ptr_deref_595_word_addrgen/root_register_ack
      -- CP-element group 128: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/ptr_deref_595_word_addrgen/root_register_req
      -- CP-element group 128: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/ptr_deref_595_word_addrgen/$exit
      -- CP-element group 128: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/ptr_deref_595_word_addrgen/$entry
      -- CP-element group 128: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/ptr_deref_595_base_plus_offset/sum_rename_ack
      -- CP-element group 128: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/ptr_deref_595_base_plus_offset/sum_rename_req
      -- CP-element group 128: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/ptr_deref_595_base_plus_offset/$exit
      -- CP-element group 128: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/ptr_deref_595_base_plus_offset/$entry
      -- CP-element group 128: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/ptr_deref_595_base_addr_resize/base_resize_ack
      -- CP-element group 128: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/ptr_deref_595_base_addr_resize/base_resize_req
      -- CP-element group 128: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/ptr_deref_595_base_addr_resize/$exit
      -- CP-element group 128: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/ptr_deref_595_base_addr_resize/$entry
      -- CP-element group 128: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/addr_of_459_update_completed_
      -- CP-element group 128: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/addr_of_459_complete/$exit
      -- CP-element group 128: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/addr_of_459_complete/ack
      -- 
    ack_1006_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_459_final_reg_ack_1, ack => convTranspose_CP_39_elements(128)); -- 
    -- CP-element group 129:  transition  input  output  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	366 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (6) 
      -- CP-element group 129: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_462_sample_completed_
      -- CP-element group 129: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_462_update_start_
      -- CP-element group 129: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_462_Sample/$exit
      -- CP-element group 129: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_462_Sample/ra
      -- CP-element group 129: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_462_Update/$entry
      -- CP-element group 129: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_462_Update/cr
      -- 
    ra_1015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_462_inst_ack_0, ack => convTranspose_CP_39_elements(129)); -- 
    cr_1019_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1019_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(129), ack => RPIPE_ConvTranspose_input_pipe_462_inst_req_1); -- 
    -- CP-element group 130:  fork  transition  input  output  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130: 	133 
    -- CP-element group 130:  members (9) 
      -- CP-element group 130: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_462_update_completed_
      -- CP-element group 130: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_462_Update/$exit
      -- CP-element group 130: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_462_Update/ca
      -- CP-element group 130: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_466_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_466_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_466_Sample/rr
      -- CP-element group 130: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_475_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_475_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_475_Sample/rr
      -- 
    ca_1020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_462_inst_ack_1, ack => convTranspose_CP_39_elements(130)); -- 
    rr_1028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(130), ack => type_cast_466_inst_req_0); -- 
    rr_1042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(130), ack => RPIPE_ConvTranspose_input_pipe_475_inst_req_0); -- 
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_466_sample_completed_
      -- CP-element group 131: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_466_Sample/$exit
      -- CP-element group 131: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_466_Sample/ra
      -- 
    ra_1029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_466_inst_ack_0, ack => convTranspose_CP_39_elements(131)); -- 
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	366 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	161 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_466_update_completed_
      -- CP-element group 132: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_466_Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_466_Update/ca
      -- 
    ca_1034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_466_inst_ack_1, ack => convTranspose_CP_39_elements(132)); -- 
    -- CP-element group 133:  transition  input  output  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	130 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133:  members (6) 
      -- CP-element group 133: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_475_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_475_update_start_
      -- CP-element group 133: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_475_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_475_Sample/ra
      -- CP-element group 133: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_475_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_475_Update/cr
      -- 
    ra_1043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_475_inst_ack_0, ack => convTranspose_CP_39_elements(133)); -- 
    cr_1047_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1047_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(133), ack => RPIPE_ConvTranspose_input_pipe_475_inst_req_1); -- 
    -- CP-element group 134:  fork  transition  input  output  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134: 	137 
    -- CP-element group 134:  members (9) 
      -- CP-element group 134: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_475_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_475_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_475_Update/ca
      -- CP-element group 134: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_479_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_479_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_479_Sample/rr
      -- CP-element group 134: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_493_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_493_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_493_Sample/rr
      -- 
    ca_1048_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_475_inst_ack_1, ack => convTranspose_CP_39_elements(134)); -- 
    rr_1070_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1070_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(134), ack => RPIPE_ConvTranspose_input_pipe_493_inst_req_0); -- 
    rr_1056_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1056_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(134), ack => type_cast_479_inst_req_0); -- 
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	134 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_479_sample_completed_
      -- CP-element group 135: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_479_Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_479_Sample/ra
      -- 
    ra_1057_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_479_inst_ack_0, ack => convTranspose_CP_39_elements(135)); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	366 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	161 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_479_update_completed_
      -- CP-element group 136: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_479_Update/$exit
      -- CP-element group 136: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_479_Update/ca
      -- 
    ca_1062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_479_inst_ack_1, ack => convTranspose_CP_39_elements(136)); -- 
    -- CP-element group 137:  transition  input  output  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	134 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137:  members (6) 
      -- CP-element group 137: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_493_sample_completed_
      -- CP-element group 137: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_493_update_start_
      -- CP-element group 137: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_493_Sample/$exit
      -- CP-element group 137: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_493_Sample/ra
      -- CP-element group 137: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_493_Update/$entry
      -- CP-element group 137: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_493_Update/cr
      -- 
    ra_1071_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_493_inst_ack_0, ack => convTranspose_CP_39_elements(137)); -- 
    cr_1075_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1075_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(137), ack => RPIPE_ConvTranspose_input_pipe_493_inst_req_1); -- 
    -- CP-element group 138:  fork  transition  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	139 
    -- CP-element group 138: 	141 
    -- CP-element group 138:  members (9) 
      -- CP-element group 138: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_493_update_completed_
      -- CP-element group 138: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_493_Update/$exit
      -- CP-element group 138: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_493_Update/ca
      -- CP-element group 138: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_497_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_497_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_497_Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_511_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_511_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_511_Sample/rr
      -- 
    ca_1076_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_493_inst_ack_1, ack => convTranspose_CP_39_elements(138)); -- 
    rr_1084_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1084_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(138), ack => type_cast_497_inst_req_0); -- 
    rr_1098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(138), ack => RPIPE_ConvTranspose_input_pipe_511_inst_req_0); -- 
    -- CP-element group 139:  transition  input  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	138 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_497_sample_completed_
      -- CP-element group 139: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_497_Sample/$exit
      -- CP-element group 139: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_497_Sample/ra
      -- 
    ra_1085_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_497_inst_ack_0, ack => convTranspose_CP_39_elements(139)); -- 
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	366 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	161 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_497_update_completed_
      -- CP-element group 140: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_497_Update/$exit
      -- CP-element group 140: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_497_Update/ca
      -- 
    ca_1090_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_497_inst_ack_1, ack => convTranspose_CP_39_elements(140)); -- 
    -- CP-element group 141:  transition  input  output  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	138 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	142 
    -- CP-element group 141:  members (6) 
      -- CP-element group 141: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_511_Update/cr
      -- CP-element group 141: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_511_Update/$entry
      -- CP-element group 141: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_511_sample_completed_
      -- CP-element group 141: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_511_update_start_
      -- CP-element group 141: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_511_Sample/$exit
      -- CP-element group 141: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_511_Sample/ra
      -- 
    ra_1099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_511_inst_ack_0, ack => convTranspose_CP_39_elements(141)); -- 
    cr_1103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(141), ack => RPIPE_ConvTranspose_input_pipe_511_inst_req_1); -- 
    -- CP-element group 142:  fork  transition  input  output  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	141 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	143 
    -- CP-element group 142: 	145 
    -- CP-element group 142:  members (9) 
      -- CP-element group 142: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_529_Sample/rr
      -- CP-element group 142: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_529_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_529_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_515_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_515_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_511_Update/ca
      -- CP-element group 142: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_511_Update/$exit
      -- CP-element group 142: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_515_Sample/rr
      -- CP-element group 142: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_511_update_completed_
      -- 
    ca_1104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_511_inst_ack_1, ack => convTranspose_CP_39_elements(142)); -- 
    rr_1112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(142), ack => type_cast_515_inst_req_0); -- 
    rr_1126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(142), ack => RPIPE_ConvTranspose_input_pipe_529_inst_req_0); -- 
    -- CP-element group 143:  transition  input  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	142 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_515_Sample/$exit
      -- CP-element group 143: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_515_Sample/ra
      -- CP-element group 143: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_515_sample_completed_
      -- 
    ra_1113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_515_inst_ack_0, ack => convTranspose_CP_39_elements(143)); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	366 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	161 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_515_Update/ca
      -- CP-element group 144: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_515_Update/$exit
      -- CP-element group 144: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_515_update_completed_
      -- 
    ca_1118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_515_inst_ack_1, ack => convTranspose_CP_39_elements(144)); -- 
    -- CP-element group 145:  transition  input  output  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	142 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145:  members (6) 
      -- CP-element group 145: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_529_Update/$entry
      -- CP-element group 145: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_529_Sample/ra
      -- CP-element group 145: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_529_Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_529_update_start_
      -- CP-element group 145: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_529_sample_completed_
      -- CP-element group 145: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_529_Update/cr
      -- 
    ra_1127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_529_inst_ack_0, ack => convTranspose_CP_39_elements(145)); -- 
    cr_1131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(145), ack => RPIPE_ConvTranspose_input_pipe_529_inst_req_1); -- 
    -- CP-element group 146:  fork  transition  input  output  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	145 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	147 
    -- CP-element group 146: 	149 
    -- CP-element group 146:  members (9) 
      -- CP-element group 146: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_529_update_completed_
      -- CP-element group 146: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_547_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_547_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_547_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_533_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_533_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_533_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_529_Update/ca
      -- CP-element group 146: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_529_Update/$exit
      -- 
    ca_1132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_529_inst_ack_1, ack => convTranspose_CP_39_elements(146)); -- 
    rr_1140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(146), ack => type_cast_533_inst_req_0); -- 
    rr_1154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(146), ack => RPIPE_ConvTranspose_input_pipe_547_inst_req_0); -- 
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	146 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_533_Sample/ra
      -- CP-element group 147: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_533_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_533_sample_completed_
      -- 
    ra_1141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_533_inst_ack_0, ack => convTranspose_CP_39_elements(147)); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	366 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	161 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_533_Update/ca
      -- CP-element group 148: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_533_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_533_update_completed_
      -- 
    ca_1146_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_533_inst_ack_1, ack => convTranspose_CP_39_elements(148)); -- 
    -- CP-element group 149:  transition  input  output  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	146 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	150 
    -- CP-element group 149:  members (6) 
      -- CP-element group 149: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_547_Update/cr
      -- CP-element group 149: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_547_Update/$entry
      -- CP-element group 149: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_547_Sample/ra
      -- CP-element group 149: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_547_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_547_update_start_
      -- CP-element group 149: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_547_sample_completed_
      -- 
    ra_1155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_547_inst_ack_0, ack => convTranspose_CP_39_elements(149)); -- 
    cr_1159_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1159_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(149), ack => RPIPE_ConvTranspose_input_pipe_547_inst_req_1); -- 
    -- CP-element group 150:  fork  transition  input  output  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	149 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	151 
    -- CP-element group 150: 	153 
    -- CP-element group 150:  members (9) 
      -- CP-element group 150: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_565_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_565_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_565_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_551_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_551_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_551_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_547_Update/ca
      -- CP-element group 150: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_547_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_547_update_completed_
      -- 
    ca_1160_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_547_inst_ack_1, ack => convTranspose_CP_39_elements(150)); -- 
    rr_1168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(150), ack => type_cast_551_inst_req_0); -- 
    rr_1182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(150), ack => RPIPE_ConvTranspose_input_pipe_565_inst_req_0); -- 
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	150 
    -- CP-element group 151: successors 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_551_Sample/ra
      -- CP-element group 151: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_551_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_551_sample_completed_
      -- 
    ra_1169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_551_inst_ack_0, ack => convTranspose_CP_39_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	366 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	161 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_551_Update/ca
      -- CP-element group 152: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_551_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_551_update_completed_
      -- 
    ca_1174_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_551_inst_ack_1, ack => convTranspose_CP_39_elements(152)); -- 
    -- CP-element group 153:  transition  input  output  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	150 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153:  members (6) 
      -- CP-element group 153: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_565_Update/cr
      -- CP-element group 153: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_565_Update/$entry
      -- CP-element group 153: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_565_Sample/ra
      -- CP-element group 153: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_565_Sample/$exit
      -- CP-element group 153: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_565_update_start_
      -- CP-element group 153: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_565_sample_completed_
      -- 
    ra_1183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_565_inst_ack_0, ack => convTranspose_CP_39_elements(153)); -- 
    cr_1187_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1187_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(153), ack => RPIPE_ConvTranspose_input_pipe_565_inst_req_1); -- 
    -- CP-element group 154:  fork  transition  input  output  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154: 	157 
    -- CP-element group 154:  members (9) 
      -- CP-element group 154: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_569_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_583_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_565_Update/ca
      -- CP-element group 154: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_569_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_569_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_565_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_565_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_583_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_583_Sample/$entry
      -- 
    ca_1188_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_565_inst_ack_1, ack => convTranspose_CP_39_elements(154)); -- 
    rr_1196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(154), ack => type_cast_569_inst_req_0); -- 
    rr_1210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(154), ack => RPIPE_ConvTranspose_input_pipe_583_inst_req_0); -- 
    -- CP-element group 155:  transition  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_569_sample_completed_
      -- CP-element group 155: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_569_Sample/ra
      -- CP-element group 155: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_569_Sample/$exit
      -- 
    ra_1197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_569_inst_ack_0, ack => convTranspose_CP_39_elements(155)); -- 
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	366 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	161 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_569_Update/ca
      -- CP-element group 156: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_569_Update/$exit
      -- CP-element group 156: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_569_update_completed_
      -- 
    ca_1202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_569_inst_ack_1, ack => convTranspose_CP_39_elements(156)); -- 
    -- CP-element group 157:  transition  input  output  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	154 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	158 
    -- CP-element group 157:  members (6) 
      -- CP-element group 157: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_583_update_start_
      -- CP-element group 157: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_583_sample_completed_
      -- CP-element group 157: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_583_Update/cr
      -- CP-element group 157: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_583_Update/$entry
      -- CP-element group 157: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_583_Sample/ra
      -- CP-element group 157: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_583_Sample/$exit
      -- 
    ra_1211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_583_inst_ack_0, ack => convTranspose_CP_39_elements(157)); -- 
    cr_1215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(157), ack => RPIPE_ConvTranspose_input_pipe_583_inst_req_1); -- 
    -- CP-element group 158:  transition  input  output  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	157 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	159 
    -- CP-element group 158:  members (6) 
      -- CP-element group 158: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_587_Sample/rr
      -- CP-element group 158: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_587_Sample/$entry
      -- CP-element group 158: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_587_sample_start_
      -- CP-element group 158: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_583_Update/ca
      -- CP-element group 158: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_583_Update/$exit
      -- CP-element group 158: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_583_update_completed_
      -- 
    ca_1216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_583_inst_ack_1, ack => convTranspose_CP_39_elements(158)); -- 
    rr_1224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(158), ack => type_cast_587_inst_req_0); -- 
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	158 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_587_Sample/ra
      -- CP-element group 159: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_587_Sample/$exit
      -- CP-element group 159: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_587_sample_completed_
      -- 
    ra_1225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_587_inst_ack_0, ack => convTranspose_CP_39_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	366 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	161 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_587_Update/ca
      -- CP-element group 160: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_587_Update/$exit
      -- CP-element group 160: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_587_update_completed_
      -- 
    ca_1230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_587_inst_ack_1, ack => convTranspose_CP_39_elements(160)); -- 
    -- CP-element group 161:  join  transition  output  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	136 
    -- CP-element group 161: 	140 
    -- CP-element group 161: 	132 
    -- CP-element group 161: 	144 
    -- CP-element group 161: 	148 
    -- CP-element group 161: 	152 
    -- CP-element group 161: 	156 
    -- CP-element group 161: 	160 
    -- CP-element group 161: 	128 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161:  members (9) 
      -- CP-element group 161: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/ptr_deref_595_sample_start_
      -- CP-element group 161: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/ptr_deref_595_Sample/word_access_start/word_0/rr
      -- CP-element group 161: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/ptr_deref_595_Sample/word_access_start/word_0/$entry
      -- CP-element group 161: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/ptr_deref_595_Sample/word_access_start/$entry
      -- CP-element group 161: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/ptr_deref_595_Sample/ptr_deref_595_Split/split_ack
      -- CP-element group 161: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/ptr_deref_595_Sample/ptr_deref_595_Split/split_req
      -- CP-element group 161: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/ptr_deref_595_Sample/ptr_deref_595_Split/$exit
      -- CP-element group 161: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/ptr_deref_595_Sample/ptr_deref_595_Split/$entry
      -- CP-element group 161: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/ptr_deref_595_Sample/$entry
      -- 
    rr_1268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(161), ack => ptr_deref_595_store_0_req_0); -- 
    convTranspose_cp_element_group_161: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_161"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(136) & convTranspose_CP_39_elements(140) & convTranspose_CP_39_elements(132) & convTranspose_CP_39_elements(144) & convTranspose_CP_39_elements(148) & convTranspose_CP_39_elements(152) & convTranspose_CP_39_elements(156) & convTranspose_CP_39_elements(160) & convTranspose_CP_39_elements(128);
      gj_convTranspose_cp_element_group_161 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(161), clk => clk, reset => reset); --
    end block;
    -- CP-element group 162:  transition  input  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	161 
    -- CP-element group 162: successors 
    -- CP-element group 162:  members (5) 
      -- CP-element group 162: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/ptr_deref_595_sample_completed_
      -- CP-element group 162: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/ptr_deref_595_Sample/word_access_start/word_0/ra
      -- CP-element group 162: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/ptr_deref_595_Sample/word_access_start/word_0/$exit
      -- CP-element group 162: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/ptr_deref_595_Sample/word_access_start/$exit
      -- CP-element group 162: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/ptr_deref_595_Sample/$exit
      -- 
    ra_1269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_595_store_0_ack_0, ack => convTranspose_CP_39_elements(162)); -- 
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	366 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	164 
    -- CP-element group 163:  members (5) 
      -- CP-element group 163: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/ptr_deref_595_update_completed_
      -- CP-element group 163: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/ptr_deref_595_Update/$exit
      -- CP-element group 163: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/ptr_deref_595_Update/word_access_complete/word_0/ca
      -- CP-element group 163: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/ptr_deref_595_Update/word_access_complete/word_0/$exit
      -- CP-element group 163: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/ptr_deref_595_Update/word_access_complete/$exit
      -- 
    ca_1280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_595_store_0_ack_1, ack => convTranspose_CP_39_elements(163)); -- 
    -- CP-element group 164:  branch  join  transition  place  output  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	163 
    -- CP-element group 164: 	125 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	165 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (10) 
      -- CP-element group 164: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608__exit__
      -- CP-element group 164: 	 branch_block_stmt_26/if_stmt_609__entry__
      -- CP-element group 164: 	 branch_block_stmt_26/if_stmt_609_else_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_26/if_stmt_609_if_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_26/R_exitcond3_610_place
      -- CP-element group 164: 	 branch_block_stmt_26/if_stmt_609_eval_test/branch_req
      -- CP-element group 164: 	 branch_block_stmt_26/if_stmt_609_eval_test/$exit
      -- CP-element group 164: 	 branch_block_stmt_26/if_stmt_609_eval_test/$entry
      -- CP-element group 164: 	 branch_block_stmt_26/if_stmt_609_dead_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/$exit
      -- 
    branch_req_1288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(164), ack => if_stmt_609_branch_req_0); -- 
    convTranspose_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(163) & convTranspose_CP_39_elements(125);
      gj_convTranspose_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  merge  transition  place  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	164 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	360 
    -- CP-element group 165:  members (13) 
      -- CP-element group 165: 	 branch_block_stmt_26/merge_stmt_393__exit__
      -- CP-element group 165: 	 branch_block_stmt_26/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader
      -- CP-element group 165: 	 branch_block_stmt_26/if_stmt_609_if_link/if_choice_transition
      -- CP-element group 165: 	 branch_block_stmt_26/if_stmt_609_if_link/$exit
      -- CP-element group 165: 	 branch_block_stmt_26/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit
      -- CP-element group 165: 	 branch_block_stmt_26/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit_PhiReq/$entry
      -- CP-element group 165: 	 branch_block_stmt_26/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit_PhiReq/$exit
      -- CP-element group 165: 	 branch_block_stmt_26/merge_stmt_393_PhiReqMerge
      -- CP-element group 165: 	 branch_block_stmt_26/merge_stmt_393_PhiAck/$entry
      -- CP-element group 165: 	 branch_block_stmt_26/merge_stmt_393_PhiAck/$exit
      -- CP-element group 165: 	 branch_block_stmt_26/merge_stmt_393_PhiAck/dummy
      -- CP-element group 165: 	 branch_block_stmt_26/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader_PhiReq/$entry
      -- CP-element group 165: 	 branch_block_stmt_26/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader_PhiReq/$exit
      -- 
    if_choice_transition_1293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_609_branch_ack_1, ack => convTranspose_CP_39_elements(165)); -- 
    -- CP-element group 166:  fork  transition  place  input  output  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	362 
    -- CP-element group 166: 	363 
    -- CP-element group 166:  members (12) 
      -- CP-element group 166: 	 branch_block_stmt_26/if_stmt_609_else_link/else_choice_transition
      -- CP-element group 166: 	 branch_block_stmt_26/if_stmt_609_else_link/$exit
      -- CP-element group 166: 	 branch_block_stmt_26/forx_xbody_forx_xbody
      -- CP-element group 166: 	 branch_block_stmt_26/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 166: 	 branch_block_stmt_26/forx_xbody_forx_xbody_PhiReq/phi_stmt_446/$entry
      -- CP-element group 166: 	 branch_block_stmt_26/forx_xbody_forx_xbody_PhiReq/phi_stmt_446/phi_stmt_446_sources/$entry
      -- CP-element group 166: 	 branch_block_stmt_26/forx_xbody_forx_xbody_PhiReq/phi_stmt_446/phi_stmt_446_sources/type_cast_452/$entry
      -- CP-element group 166: 	 branch_block_stmt_26/forx_xbody_forx_xbody_PhiReq/phi_stmt_446/phi_stmt_446_sources/type_cast_452/SplitProtocol/$entry
      -- CP-element group 166: 	 branch_block_stmt_26/forx_xbody_forx_xbody_PhiReq/phi_stmt_446/phi_stmt_446_sources/type_cast_452/SplitProtocol/Sample/$entry
      -- CP-element group 166: 	 branch_block_stmt_26/forx_xbody_forx_xbody_PhiReq/phi_stmt_446/phi_stmt_446_sources/type_cast_452/SplitProtocol/Sample/rr
      -- CP-element group 166: 	 branch_block_stmt_26/forx_xbody_forx_xbody_PhiReq/phi_stmt_446/phi_stmt_446_sources/type_cast_452/SplitProtocol/Update/$entry
      -- CP-element group 166: 	 branch_block_stmt_26/forx_xbody_forx_xbody_PhiReq/phi_stmt_446/phi_stmt_446_sources/type_cast_452/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1297_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_609_branch_ack_0, ack => convTranspose_CP_39_elements(166)); -- 
    rr_2802_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2802_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(166), ack => type_cast_452_inst_req_0); -- 
    cr_2807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(166), ack => type_cast_452_inst_req_1); -- 
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	121 
    -- CP-element group 167: successors 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_26/assign_stmt_621_to_assign_stmt_650/type_cast_636_Sample/ra
      -- CP-element group 167: 	 branch_block_stmt_26/assign_stmt_621_to_assign_stmt_650/type_cast_636_Sample/$exit
      -- CP-element group 167: 	 branch_block_stmt_26/assign_stmt_621_to_assign_stmt_650/type_cast_636_sample_completed_
      -- 
    ra_1311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_636_inst_ack_0, ack => convTranspose_CP_39_elements(167)); -- 
    -- CP-element group 168:  transition  place  input  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	121 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	367 
    -- CP-element group 168:  members (9) 
      -- CP-element group 168: 	 branch_block_stmt_26/assign_stmt_621_to_assign_stmt_650__exit__
      -- CP-element group 168: 	 branch_block_stmt_26/bbx_xnph454_forx_xbody196
      -- CP-element group 168: 	 branch_block_stmt_26/assign_stmt_621_to_assign_stmt_650/type_cast_636_Update/ca
      -- CP-element group 168: 	 branch_block_stmt_26/assign_stmt_621_to_assign_stmt_650/type_cast_636_Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_26/assign_stmt_621_to_assign_stmt_650/type_cast_636_update_completed_
      -- CP-element group 168: 	 branch_block_stmt_26/assign_stmt_621_to_assign_stmt_650/$exit
      -- CP-element group 168: 	 branch_block_stmt_26/bbx_xnph454_forx_xbody196_PhiReq/$entry
      -- CP-element group 168: 	 branch_block_stmt_26/bbx_xnph454_forx_xbody196_PhiReq/phi_stmt_653/$entry
      -- CP-element group 168: 	 branch_block_stmt_26/bbx_xnph454_forx_xbody196_PhiReq/phi_stmt_653/phi_stmt_653_sources/$entry
      -- 
    ca_1316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_636_inst_ack_1, ack => convTranspose_CP_39_elements(168)); -- 
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	372 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	208 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/array_obj_ref_665_final_index_sum_regn_Sample/ack
      -- CP-element group 169: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/array_obj_ref_665_final_index_sum_regn_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/array_obj_ref_665_final_index_sum_regn_sample_complete
      -- 
    ack_1345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_665_index_offset_ack_0, ack => convTranspose_CP_39_elements(169)); -- 
    -- CP-element group 170:  transition  input  output  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	372 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	171 
    -- CP-element group 170:  members (11) 
      -- CP-element group 170: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/array_obj_ref_665_offset_calculated
      -- CP-element group 170: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/addr_of_666_request/req
      -- CP-element group 170: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/array_obj_ref_665_root_address_calculated
      -- CP-element group 170: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/addr_of_666_request/$entry
      -- CP-element group 170: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/array_obj_ref_665_base_plus_offset/sum_rename_ack
      -- CP-element group 170: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/addr_of_666_sample_start_
      -- CP-element group 170: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/array_obj_ref_665_base_plus_offset/sum_rename_req
      -- CP-element group 170: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/array_obj_ref_665_base_plus_offset/$exit
      -- CP-element group 170: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/array_obj_ref_665_base_plus_offset/$entry
      -- CP-element group 170: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/array_obj_ref_665_final_index_sum_regn_Update/ack
      -- CP-element group 170: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/array_obj_ref_665_final_index_sum_regn_Update/$exit
      -- 
    ack_1350_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_665_index_offset_ack_1, ack => convTranspose_CP_39_elements(170)); -- 
    req_1359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(170), ack => addr_of_666_final_reg_req_0); -- 
    -- CP-element group 171:  transition  input  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	170 
    -- CP-element group 171: successors 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/addr_of_666_request/$exit
      -- CP-element group 171: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/addr_of_666_sample_completed_
      -- CP-element group 171: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/addr_of_666_request/ack
      -- 
    ack_1360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_666_final_reg_ack_0, ack => convTranspose_CP_39_elements(171)); -- 
    -- CP-element group 172:  fork  transition  input  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	372 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	205 
    -- CP-element group 172:  members (19) 
      -- CP-element group 172: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/addr_of_666_update_completed_
      -- CP-element group 172: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/addr_of_666_complete/ack
      -- CP-element group 172: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/addr_of_666_complete/$exit
      -- CP-element group 172: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/ptr_deref_802_base_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/ptr_deref_802_word_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/ptr_deref_802_root_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/ptr_deref_802_base_address_resized
      -- CP-element group 172: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/ptr_deref_802_base_addr_resize/$entry
      -- CP-element group 172: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/ptr_deref_802_base_addr_resize/$exit
      -- CP-element group 172: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/ptr_deref_802_base_addr_resize/base_resize_req
      -- CP-element group 172: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/ptr_deref_802_base_addr_resize/base_resize_ack
      -- CP-element group 172: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/ptr_deref_802_base_plus_offset/$entry
      -- CP-element group 172: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/ptr_deref_802_base_plus_offset/$exit
      -- CP-element group 172: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/ptr_deref_802_base_plus_offset/sum_rename_req
      -- CP-element group 172: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/ptr_deref_802_base_plus_offset/sum_rename_ack
      -- CP-element group 172: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/ptr_deref_802_word_addrgen/$entry
      -- CP-element group 172: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/ptr_deref_802_word_addrgen/$exit
      -- CP-element group 172: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/ptr_deref_802_word_addrgen/root_register_req
      -- CP-element group 172: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/ptr_deref_802_word_addrgen/root_register_ack
      -- 
    ack_1365_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_666_final_reg_ack_1, ack => convTranspose_CP_39_elements(172)); -- 
    -- CP-element group 173:  transition  input  output  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	372 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	174 
    -- CP-element group 173:  members (6) 
      -- CP-element group 173: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_669_update_start_
      -- CP-element group 173: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_669_sample_completed_
      -- CP-element group 173: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_669_Update/cr
      -- CP-element group 173: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_669_Update/$entry
      -- CP-element group 173: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_669_Sample/ra
      -- CP-element group 173: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_669_Sample/$exit
      -- 
    ra_1374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_669_inst_ack_0, ack => convTranspose_CP_39_elements(173)); -- 
    cr_1378_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1378_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(173), ack => RPIPE_ConvTranspose_input_pipe_669_inst_req_1); -- 
    -- CP-element group 174:  fork  transition  input  output  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	173 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	175 
    -- CP-element group 174: 	177 
    -- CP-element group 174:  members (9) 
      -- CP-element group 174: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_673_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_669_update_completed_
      -- CP-element group 174: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_669_Update/ca
      -- CP-element group 174: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_673_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_669_Update/$exit
      -- CP-element group 174: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_682_Sample/rr
      -- CP-element group 174: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_682_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_682_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_673_Sample/rr
      -- 
    ca_1379_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_669_inst_ack_1, ack => convTranspose_CP_39_elements(174)); -- 
    rr_1387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(174), ack => type_cast_673_inst_req_0); -- 
    rr_1401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(174), ack => RPIPE_ConvTranspose_input_pipe_682_inst_req_0); -- 
    -- CP-element group 175:  transition  input  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	174 
    -- CP-element group 175: successors 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_673_sample_completed_
      -- CP-element group 175: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_673_Sample/ra
      -- CP-element group 175: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_673_Sample/$exit
      -- 
    ra_1388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_673_inst_ack_0, ack => convTranspose_CP_39_elements(175)); -- 
    -- CP-element group 176:  transition  input  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	372 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	205 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_673_update_completed_
      -- CP-element group 176: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_673_Update/ca
      -- CP-element group 176: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_673_Update/$exit
      -- 
    ca_1393_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_673_inst_ack_1, ack => convTranspose_CP_39_elements(176)); -- 
    -- CP-element group 177:  transition  input  output  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	174 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	178 
    -- CP-element group 177:  members (6) 
      -- CP-element group 177: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_682_Update/cr
      -- CP-element group 177: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_682_Update/$entry
      -- CP-element group 177: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_682_Sample/ra
      -- CP-element group 177: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_682_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_682_update_start_
      -- CP-element group 177: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_682_sample_completed_
      -- 
    ra_1402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_682_inst_ack_0, ack => convTranspose_CP_39_elements(177)); -- 
    cr_1406_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1406_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(177), ack => RPIPE_ConvTranspose_input_pipe_682_inst_req_1); -- 
    -- CP-element group 178:  fork  transition  input  output  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	177 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178: 	181 
    -- CP-element group 178:  members (9) 
      -- CP-element group 178: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_686_sample_start_
      -- CP-element group 178: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_686_Sample/$entry
      -- CP-element group 178: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_700_sample_start_
      -- CP-element group 178: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_682_Update/ca
      -- CP-element group 178: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_682_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_686_Sample/rr
      -- CP-element group 178: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_682_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_700_Sample/rr
      -- CP-element group 178: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_700_Sample/$entry
      -- 
    ca_1407_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_682_inst_ack_1, ack => convTranspose_CP_39_elements(178)); -- 
    rr_1415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(178), ack => type_cast_686_inst_req_0); -- 
    rr_1429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(178), ack => RPIPE_ConvTranspose_input_pipe_700_inst_req_0); -- 
    -- CP-element group 179:  transition  input  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	178 
    -- CP-element group 179: successors 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_686_sample_completed_
      -- CP-element group 179: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_686_Sample/ra
      -- CP-element group 179: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_686_Sample/$exit
      -- 
    ra_1416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_686_inst_ack_0, ack => convTranspose_CP_39_elements(179)); -- 
    -- CP-element group 180:  transition  input  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	372 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	205 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_686_Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_686_update_completed_
      -- CP-element group 180: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_686_Update/ca
      -- 
    ca_1421_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_686_inst_ack_1, ack => convTranspose_CP_39_elements(180)); -- 
    -- CP-element group 181:  transition  input  output  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	178 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	182 
    -- CP-element group 181:  members (6) 
      -- CP-element group 181: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_700_sample_completed_
      -- CP-element group 181: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_700_Update/cr
      -- CP-element group 181: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_700_Update/$entry
      -- CP-element group 181: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_700_Sample/ra
      -- CP-element group 181: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_700_Sample/$exit
      -- CP-element group 181: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_700_update_start_
      -- 
    ra_1430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_700_inst_ack_0, ack => convTranspose_CP_39_elements(181)); -- 
    cr_1434_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1434_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(181), ack => RPIPE_ConvTranspose_input_pipe_700_inst_req_1); -- 
    -- CP-element group 182:  fork  transition  input  output  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	181 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	183 
    -- CP-element group 182: 	185 
    -- CP-element group 182:  members (9) 
      -- CP-element group 182: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_718_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_704_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_718_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_718_Sample/rr
      -- CP-element group 182: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_700_Update/ca
      -- CP-element group 182: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_704_Sample/rr
      -- CP-element group 182: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_700_Update/$exit
      -- CP-element group 182: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_704_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_700_update_completed_
      -- 
    ca_1435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_700_inst_ack_1, ack => convTranspose_CP_39_elements(182)); -- 
    rr_1443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(182), ack => type_cast_704_inst_req_0); -- 
    rr_1457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(182), ack => RPIPE_ConvTranspose_input_pipe_718_inst_req_0); -- 
    -- CP-element group 183:  transition  input  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	182 
    -- CP-element group 183: successors 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_704_sample_completed_
      -- CP-element group 183: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_704_Sample/ra
      -- CP-element group 183: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_704_Sample/$exit
      -- 
    ra_1444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_704_inst_ack_0, ack => convTranspose_CP_39_elements(183)); -- 
    -- CP-element group 184:  transition  input  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	372 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	205 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_704_Update/ca
      -- CP-element group 184: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_704_Update/$exit
      -- CP-element group 184: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_704_update_completed_
      -- 
    ca_1449_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_704_inst_ack_1, ack => convTranspose_CP_39_elements(184)); -- 
    -- CP-element group 185:  transition  input  output  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	182 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	186 
    -- CP-element group 185:  members (6) 
      -- CP-element group 185: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_718_Sample/$exit
      -- CP-element group 185: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_718_Update/$entry
      -- CP-element group 185: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_718_update_start_
      -- CP-element group 185: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_718_Update/cr
      -- CP-element group 185: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_718_sample_completed_
      -- CP-element group 185: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_718_Sample/ra
      -- 
    ra_1458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_718_inst_ack_0, ack => convTranspose_CP_39_elements(185)); -- 
    cr_1462_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1462_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(185), ack => RPIPE_ConvTranspose_input_pipe_718_inst_req_1); -- 
    -- CP-element group 186:  fork  transition  input  output  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	185 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186: 	189 
    -- CP-element group 186:  members (9) 
      -- CP-element group 186: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_718_update_completed_
      -- CP-element group 186: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_718_Update/$exit
      -- CP-element group 186: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_722_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_718_Update/ca
      -- CP-element group 186: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_722_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_722_Sample/rr
      -- CP-element group 186: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_736_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_736_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_736_Sample/rr
      -- 
    ca_1463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_718_inst_ack_1, ack => convTranspose_CP_39_elements(186)); -- 
    rr_1471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(186), ack => type_cast_722_inst_req_0); -- 
    rr_1485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(186), ack => RPIPE_ConvTranspose_input_pipe_736_inst_req_0); -- 
    -- CP-element group 187:  transition  input  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_722_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_722_Sample/$exit
      -- CP-element group 187: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_722_Sample/ra
      -- 
    ra_1472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_722_inst_ack_0, ack => convTranspose_CP_39_elements(187)); -- 
    -- CP-element group 188:  transition  input  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	372 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	205 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_722_update_completed_
      -- CP-element group 188: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_722_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_722_Update/ca
      -- 
    ca_1477_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_722_inst_ack_1, ack => convTranspose_CP_39_elements(188)); -- 
    -- CP-element group 189:  transition  input  output  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	186 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	190 
    -- CP-element group 189:  members (6) 
      -- CP-element group 189: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_736_sample_completed_
      -- CP-element group 189: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_736_update_start_
      -- CP-element group 189: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_736_Sample/$exit
      -- CP-element group 189: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_736_Sample/ra
      -- CP-element group 189: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_736_Update/$entry
      -- CP-element group 189: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_736_Update/cr
      -- 
    ra_1486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_736_inst_ack_0, ack => convTranspose_CP_39_elements(189)); -- 
    cr_1490_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1490_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(189), ack => RPIPE_ConvTranspose_input_pipe_736_inst_req_1); -- 
    -- CP-element group 190:  fork  transition  input  output  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	189 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	191 
    -- CP-element group 190: 	193 
    -- CP-element group 190:  members (9) 
      -- CP-element group 190: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_736_update_completed_
      -- CP-element group 190: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_736_Update/$exit
      -- CP-element group 190: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_736_Update/ca
      -- CP-element group 190: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_740_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_740_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_740_Sample/rr
      -- CP-element group 190: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_754_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_754_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_754_Sample/rr
      -- 
    ca_1491_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_736_inst_ack_1, ack => convTranspose_CP_39_elements(190)); -- 
    rr_1499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(190), ack => type_cast_740_inst_req_0); -- 
    rr_1513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(190), ack => RPIPE_ConvTranspose_input_pipe_754_inst_req_0); -- 
    -- CP-element group 191:  transition  input  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	190 
    -- CP-element group 191: successors 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_740_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_740_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_740_Sample/ra
      -- 
    ra_1500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_740_inst_ack_0, ack => convTranspose_CP_39_elements(191)); -- 
    -- CP-element group 192:  transition  input  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	372 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	205 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_740_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_740_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_740_Update/ca
      -- 
    ca_1505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_740_inst_ack_1, ack => convTranspose_CP_39_elements(192)); -- 
    -- CP-element group 193:  transition  input  output  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	190 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	194 
    -- CP-element group 193:  members (6) 
      -- CP-element group 193: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_754_sample_completed_
      -- CP-element group 193: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_754_update_start_
      -- CP-element group 193: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_754_Sample/$exit
      -- CP-element group 193: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_754_Sample/ra
      -- CP-element group 193: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_754_Update/$entry
      -- CP-element group 193: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_754_Update/cr
      -- 
    ra_1514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_754_inst_ack_0, ack => convTranspose_CP_39_elements(193)); -- 
    cr_1518_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1518_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(193), ack => RPIPE_ConvTranspose_input_pipe_754_inst_req_1); -- 
    -- CP-element group 194:  fork  transition  input  output  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	193 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194: 	197 
    -- CP-element group 194:  members (9) 
      -- CP-element group 194: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_754_update_completed_
      -- CP-element group 194: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_754_Update/$exit
      -- CP-element group 194: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_754_Update/ca
      -- CP-element group 194: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_758_sample_start_
      -- CP-element group 194: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_758_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_758_Sample/rr
      -- CP-element group 194: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_772_sample_start_
      -- CP-element group 194: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_772_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_772_Sample/rr
      -- 
    ca_1519_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_754_inst_ack_1, ack => convTranspose_CP_39_elements(194)); -- 
    rr_1527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(194), ack => type_cast_758_inst_req_0); -- 
    rr_1541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(194), ack => RPIPE_ConvTranspose_input_pipe_772_inst_req_0); -- 
    -- CP-element group 195:  transition  input  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_758_sample_completed_
      -- CP-element group 195: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_758_Sample/$exit
      -- CP-element group 195: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_758_Sample/ra
      -- 
    ra_1528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_758_inst_ack_0, ack => convTranspose_CP_39_elements(195)); -- 
    -- CP-element group 196:  transition  input  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	372 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	205 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_758_update_completed_
      -- CP-element group 196: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_758_Update/$exit
      -- CP-element group 196: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_758_Update/ca
      -- 
    ca_1533_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_758_inst_ack_1, ack => convTranspose_CP_39_elements(196)); -- 
    -- CP-element group 197:  transition  input  output  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	194 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	198 
    -- CP-element group 197:  members (6) 
      -- CP-element group 197: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_772_sample_completed_
      -- CP-element group 197: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_772_update_start_
      -- CP-element group 197: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_772_Sample/$exit
      -- CP-element group 197: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_772_Sample/ra
      -- CP-element group 197: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_772_Update/$entry
      -- CP-element group 197: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_772_Update/cr
      -- 
    ra_1542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_772_inst_ack_0, ack => convTranspose_CP_39_elements(197)); -- 
    cr_1546_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1546_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(197), ack => RPIPE_ConvTranspose_input_pipe_772_inst_req_1); -- 
    -- CP-element group 198:  fork  transition  input  output  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	197 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	199 
    -- CP-element group 198: 	201 
    -- CP-element group 198:  members (9) 
      -- CP-element group 198: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_772_update_completed_
      -- CP-element group 198: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_772_Update/$exit
      -- CP-element group 198: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_772_Update/ca
      -- CP-element group 198: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_776_sample_start_
      -- CP-element group 198: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_776_Sample/$entry
      -- CP-element group 198: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_776_Sample/rr
      -- CP-element group 198: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_790_sample_start_
      -- CP-element group 198: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_790_Sample/$entry
      -- CP-element group 198: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_790_Sample/rr
      -- 
    ca_1547_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_772_inst_ack_1, ack => convTranspose_CP_39_elements(198)); -- 
    rr_1555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(198), ack => type_cast_776_inst_req_0); -- 
    rr_1569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(198), ack => RPIPE_ConvTranspose_input_pipe_790_inst_req_0); -- 
    -- CP-element group 199:  transition  input  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	198 
    -- CP-element group 199: successors 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_776_sample_completed_
      -- CP-element group 199: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_776_Sample/$exit
      -- CP-element group 199: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_776_Sample/ra
      -- 
    ra_1556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_776_inst_ack_0, ack => convTranspose_CP_39_elements(199)); -- 
    -- CP-element group 200:  transition  input  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	372 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	205 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_776_update_completed_
      -- CP-element group 200: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_776_Update/$exit
      -- CP-element group 200: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_776_Update/ca
      -- 
    ca_1561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_776_inst_ack_1, ack => convTranspose_CP_39_elements(200)); -- 
    -- CP-element group 201:  transition  input  output  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	198 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201:  members (6) 
      -- CP-element group 201: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_790_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_790_update_start_
      -- CP-element group 201: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_790_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_790_Sample/ra
      -- CP-element group 201: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_790_Update/$entry
      -- CP-element group 201: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_790_Update/cr
      -- 
    ra_1570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_790_inst_ack_0, ack => convTranspose_CP_39_elements(201)); -- 
    cr_1574_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1574_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(201), ack => RPIPE_ConvTranspose_input_pipe_790_inst_req_1); -- 
    -- CP-element group 202:  transition  input  output  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	201 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202:  members (6) 
      -- CP-element group 202: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_790_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_790_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_790_Update/ca
      -- CP-element group 202: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_794_sample_start_
      -- CP-element group 202: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_794_Sample/$entry
      -- CP-element group 202: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_794_Sample/rr
      -- 
    ca_1575_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_790_inst_ack_1, ack => convTranspose_CP_39_elements(202)); -- 
    rr_1583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(202), ack => type_cast_794_inst_req_0); -- 
    -- CP-element group 203:  transition  input  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	202 
    -- CP-element group 203: successors 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_794_sample_completed_
      -- CP-element group 203: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_794_Sample/$exit
      -- CP-element group 203: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_794_Sample/ra
      -- 
    ra_1584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_794_inst_ack_0, ack => convTranspose_CP_39_elements(203)); -- 
    -- CP-element group 204:  transition  input  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	372 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	205 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_794_update_completed_
      -- CP-element group 204: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_794_Update/$exit
      -- CP-element group 204: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_794_Update/ca
      -- 
    ca_1589_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_794_inst_ack_1, ack => convTranspose_CP_39_elements(204)); -- 
    -- CP-element group 205:  join  transition  output  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	172 
    -- CP-element group 205: 	176 
    -- CP-element group 205: 	180 
    -- CP-element group 205: 	184 
    -- CP-element group 205: 	188 
    -- CP-element group 205: 	192 
    -- CP-element group 205: 	196 
    -- CP-element group 205: 	200 
    -- CP-element group 205: 	204 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	206 
    -- CP-element group 205:  members (9) 
      -- CP-element group 205: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/ptr_deref_802_sample_start_
      -- CP-element group 205: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/ptr_deref_802_Sample/$entry
      -- CP-element group 205: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/ptr_deref_802_Sample/ptr_deref_802_Split/$entry
      -- CP-element group 205: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/ptr_deref_802_Sample/ptr_deref_802_Split/$exit
      -- CP-element group 205: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/ptr_deref_802_Sample/ptr_deref_802_Split/split_req
      -- CP-element group 205: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/ptr_deref_802_Sample/ptr_deref_802_Split/split_ack
      -- CP-element group 205: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/ptr_deref_802_Sample/word_access_start/$entry
      -- CP-element group 205: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/ptr_deref_802_Sample/word_access_start/word_0/$entry
      -- CP-element group 205: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/ptr_deref_802_Sample/word_access_start/word_0/rr
      -- 
    rr_1627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(205), ack => ptr_deref_802_store_0_req_0); -- 
    convTranspose_cp_element_group_205: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_205"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(172) & convTranspose_CP_39_elements(176) & convTranspose_CP_39_elements(180) & convTranspose_CP_39_elements(184) & convTranspose_CP_39_elements(188) & convTranspose_CP_39_elements(192) & convTranspose_CP_39_elements(196) & convTranspose_CP_39_elements(200) & convTranspose_CP_39_elements(204);
      gj_convTranspose_cp_element_group_205 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(205), clk => clk, reset => reset); --
    end block;
    -- CP-element group 206:  transition  input  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	205 
    -- CP-element group 206: successors 
    -- CP-element group 206:  members (5) 
      -- CP-element group 206: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/ptr_deref_802_sample_completed_
      -- CP-element group 206: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/ptr_deref_802_Sample/$exit
      -- CP-element group 206: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/ptr_deref_802_Sample/word_access_start/$exit
      -- CP-element group 206: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/ptr_deref_802_Sample/word_access_start/word_0/$exit
      -- CP-element group 206: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/ptr_deref_802_Sample/word_access_start/word_0/ra
      -- 
    ra_1628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_802_store_0_ack_0, ack => convTranspose_CP_39_elements(206)); -- 
    -- CP-element group 207:  transition  input  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	372 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	208 
    -- CP-element group 207:  members (5) 
      -- CP-element group 207: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/ptr_deref_802_update_completed_
      -- CP-element group 207: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/ptr_deref_802_Update/$exit
      -- CP-element group 207: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/ptr_deref_802_Update/word_access_complete/$exit
      -- CP-element group 207: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/ptr_deref_802_Update/word_access_complete/word_0/$exit
      -- CP-element group 207: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/ptr_deref_802_Update/word_access_complete/word_0/ca
      -- 
    ca_1639_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_802_store_0_ack_1, ack => convTranspose_CP_39_elements(207)); -- 
    -- CP-element group 208:  branch  join  transition  place  output  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	169 
    -- CP-element group 208: 	207 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	209 
    -- CP-element group 208: 	210 
    -- CP-element group 208:  members (10) 
      -- CP-element group 208: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815__exit__
      -- CP-element group 208: 	 branch_block_stmt_26/if_stmt_816__entry__
      -- CP-element group 208: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/$exit
      -- CP-element group 208: 	 branch_block_stmt_26/if_stmt_816_dead_link/$entry
      -- CP-element group 208: 	 branch_block_stmt_26/if_stmt_816_eval_test/$entry
      -- CP-element group 208: 	 branch_block_stmt_26/if_stmt_816_eval_test/$exit
      -- CP-element group 208: 	 branch_block_stmt_26/if_stmt_816_eval_test/branch_req
      -- CP-element group 208: 	 branch_block_stmt_26/R_exitcond2_817_place
      -- CP-element group 208: 	 branch_block_stmt_26/if_stmt_816_if_link/$entry
      -- CP-element group 208: 	 branch_block_stmt_26/if_stmt_816_else_link/$entry
      -- 
    branch_req_1647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(208), ack => if_stmt_816_branch_req_0); -- 
    convTranspose_cp_element_group_208: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_208"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(169) & convTranspose_CP_39_elements(207);
      gj_convTranspose_cp_element_group_208 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(208), clk => clk, reset => reset); --
    end block;
    -- CP-element group 209:  merge  transition  place  input  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	208 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	373 
    -- CP-element group 209:  members (13) 
      -- CP-element group 209: 	 branch_block_stmt_26/merge_stmt_822__exit__
      -- CP-element group 209: 	 branch_block_stmt_26/forx_xend250x_xloopexit_forx_xend250
      -- CP-element group 209: 	 branch_block_stmt_26/if_stmt_816_if_link/$exit
      -- CP-element group 209: 	 branch_block_stmt_26/if_stmt_816_if_link/if_choice_transition
      -- CP-element group 209: 	 branch_block_stmt_26/forx_xbody196_forx_xend250x_xloopexit
      -- CP-element group 209: 	 branch_block_stmt_26/forx_xbody196_forx_xend250x_xloopexit_PhiReq/$entry
      -- CP-element group 209: 	 branch_block_stmt_26/forx_xbody196_forx_xend250x_xloopexit_PhiReq/$exit
      -- CP-element group 209: 	 branch_block_stmt_26/merge_stmt_822_PhiReqMerge
      -- CP-element group 209: 	 branch_block_stmt_26/merge_stmt_822_PhiAck/$entry
      -- CP-element group 209: 	 branch_block_stmt_26/merge_stmt_822_PhiAck/$exit
      -- CP-element group 209: 	 branch_block_stmt_26/merge_stmt_822_PhiAck/dummy
      -- CP-element group 209: 	 branch_block_stmt_26/forx_xend250x_xloopexit_forx_xend250_PhiReq/$entry
      -- CP-element group 209: 	 branch_block_stmt_26/forx_xend250x_xloopexit_forx_xend250_PhiReq/$exit
      -- 
    if_choice_transition_1652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_816_branch_ack_1, ack => convTranspose_CP_39_elements(209)); -- 
    -- CP-element group 210:  fork  transition  place  input  output  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	208 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	368 
    -- CP-element group 210: 	369 
    -- CP-element group 210:  members (12) 
      -- CP-element group 210: 	 branch_block_stmt_26/if_stmt_816_else_link/$exit
      -- CP-element group 210: 	 branch_block_stmt_26/if_stmt_816_else_link/else_choice_transition
      -- CP-element group 210: 	 branch_block_stmt_26/forx_xbody196_forx_xbody196
      -- CP-element group 210: 	 branch_block_stmt_26/forx_xbody196_forx_xbody196_PhiReq/$entry
      -- CP-element group 210: 	 branch_block_stmt_26/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_653/$entry
      -- CP-element group 210: 	 branch_block_stmt_26/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_653/phi_stmt_653_sources/$entry
      -- CP-element group 210: 	 branch_block_stmt_26/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_653/phi_stmt_653_sources/type_cast_659/$entry
      -- CP-element group 210: 	 branch_block_stmt_26/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_653/phi_stmt_653_sources/type_cast_659/SplitProtocol/$entry
      -- CP-element group 210: 	 branch_block_stmt_26/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_653/phi_stmt_653_sources/type_cast_659/SplitProtocol/Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_26/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_653/phi_stmt_653_sources/type_cast_659/SplitProtocol/Sample/rr
      -- CP-element group 210: 	 branch_block_stmt_26/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_653/phi_stmt_653_sources/type_cast_659/SplitProtocol/Update/$entry
      -- CP-element group 210: 	 branch_block_stmt_26/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_653/phi_stmt_653_sources/type_cast_659/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_816_branch_ack_0, ack => convTranspose_CP_39_elements(210)); -- 
    rr_2856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(210), ack => type_cast_659_inst_req_0); -- 
    cr_2861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(210), ack => type_cast_659_inst_req_1); -- 
    -- CP-element group 211:  transition  input  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	373 
    -- CP-element group 211: successors 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_26/assign_stmt_828_to_assign_stmt_852/type_cast_827_sample_completed_
      -- CP-element group 211: 	 branch_block_stmt_26/assign_stmt_828_to_assign_stmt_852/type_cast_827_Sample/$exit
      -- CP-element group 211: 	 branch_block_stmt_26/assign_stmt_828_to_assign_stmt_852/type_cast_827_Sample/ra
      -- 
    ra_1670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_827_inst_ack_0, ack => convTranspose_CP_39_elements(211)); -- 
    -- CP-element group 212:  transition  input  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	373 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	217 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_26/assign_stmt_828_to_assign_stmt_852/type_cast_827_update_completed_
      -- CP-element group 212: 	 branch_block_stmt_26/assign_stmt_828_to_assign_stmt_852/type_cast_827_Update/$exit
      -- CP-element group 212: 	 branch_block_stmt_26/assign_stmt_828_to_assign_stmt_852/type_cast_827_Update/ca
      -- 
    ca_1675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_827_inst_ack_1, ack => convTranspose_CP_39_elements(212)); -- 
    -- CP-element group 213:  transition  input  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	373 
    -- CP-element group 213: successors 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_26/assign_stmt_828_to_assign_stmt_852/type_cast_831_sample_completed_
      -- CP-element group 213: 	 branch_block_stmt_26/assign_stmt_828_to_assign_stmt_852/type_cast_831_Sample/$exit
      -- CP-element group 213: 	 branch_block_stmt_26/assign_stmt_828_to_assign_stmt_852/type_cast_831_Sample/ra
      -- 
    ra_1684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_831_inst_ack_0, ack => convTranspose_CP_39_elements(213)); -- 
    -- CP-element group 214:  transition  input  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	373 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	217 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_26/assign_stmt_828_to_assign_stmt_852/type_cast_831_update_completed_
      -- CP-element group 214: 	 branch_block_stmt_26/assign_stmt_828_to_assign_stmt_852/type_cast_831_Update/$exit
      -- CP-element group 214: 	 branch_block_stmt_26/assign_stmt_828_to_assign_stmt_852/type_cast_831_Update/ca
      -- 
    ca_1689_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_831_inst_ack_1, ack => convTranspose_CP_39_elements(214)); -- 
    -- CP-element group 215:  transition  input  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	373 
    -- CP-element group 215: successors 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_26/assign_stmt_828_to_assign_stmt_852/type_cast_835_sample_completed_
      -- CP-element group 215: 	 branch_block_stmt_26/assign_stmt_828_to_assign_stmt_852/type_cast_835_Sample/$exit
      -- CP-element group 215: 	 branch_block_stmt_26/assign_stmt_828_to_assign_stmt_852/type_cast_835_Sample/ra
      -- 
    ra_1698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_835_inst_ack_0, ack => convTranspose_CP_39_elements(215)); -- 
    -- CP-element group 216:  transition  input  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	373 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	217 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_26/assign_stmt_828_to_assign_stmt_852/type_cast_835_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_26/assign_stmt_828_to_assign_stmt_852/type_cast_835_Update/$exit
      -- CP-element group 216: 	 branch_block_stmt_26/assign_stmt_828_to_assign_stmt_852/type_cast_835_Update/ca
      -- 
    ca_1703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_835_inst_ack_1, ack => convTranspose_CP_39_elements(216)); -- 
    -- CP-element group 217:  branch  join  transition  place  output  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	212 
    -- CP-element group 217: 	214 
    -- CP-element group 217: 	216 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	218 
    -- CP-element group 217: 	219 
    -- CP-element group 217:  members (10) 
      -- CP-element group 217: 	 branch_block_stmt_26/assign_stmt_828_to_assign_stmt_852__exit__
      -- CP-element group 217: 	 branch_block_stmt_26/if_stmt_853__entry__
      -- CP-element group 217: 	 branch_block_stmt_26/assign_stmt_828_to_assign_stmt_852/$exit
      -- CP-element group 217: 	 branch_block_stmt_26/if_stmt_853_dead_link/$entry
      -- CP-element group 217: 	 branch_block_stmt_26/if_stmt_853_eval_test/$entry
      -- CP-element group 217: 	 branch_block_stmt_26/if_stmt_853_eval_test/$exit
      -- CP-element group 217: 	 branch_block_stmt_26/if_stmt_853_eval_test/branch_req
      -- CP-element group 217: 	 branch_block_stmt_26/R_cmp264448_854_place
      -- CP-element group 217: 	 branch_block_stmt_26/if_stmt_853_if_link/$entry
      -- CP-element group 217: 	 branch_block_stmt_26/if_stmt_853_else_link/$entry
      -- 
    branch_req_1711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(217), ack => if_stmt_853_branch_req_0); -- 
    convTranspose_cp_element_group_217: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_217"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(212) & convTranspose_CP_39_elements(214) & convTranspose_CP_39_elements(216);
      gj_convTranspose_cp_element_group_217 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(217), clk => clk, reset => reset); --
    end block;
    -- CP-element group 218:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	217 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	220 
    -- CP-element group 218: 	221 
    -- CP-element group 218:  members (18) 
      -- CP-element group 218: 	 branch_block_stmt_26/merge_stmt_859__exit__
      -- CP-element group 218: 	 branch_block_stmt_26/assign_stmt_865_to_assign_stmt_894__entry__
      -- CP-element group 218: 	 branch_block_stmt_26/if_stmt_853_if_link/$exit
      -- CP-element group 218: 	 branch_block_stmt_26/if_stmt_853_if_link/if_choice_transition
      -- CP-element group 218: 	 branch_block_stmt_26/forx_xend250_bbx_xnph450
      -- CP-element group 218: 	 branch_block_stmt_26/assign_stmt_865_to_assign_stmt_894/$entry
      -- CP-element group 218: 	 branch_block_stmt_26/assign_stmt_865_to_assign_stmt_894/type_cast_880_sample_start_
      -- CP-element group 218: 	 branch_block_stmt_26/assign_stmt_865_to_assign_stmt_894/type_cast_880_update_start_
      -- CP-element group 218: 	 branch_block_stmt_26/assign_stmt_865_to_assign_stmt_894/type_cast_880_Sample/$entry
      -- CP-element group 218: 	 branch_block_stmt_26/assign_stmt_865_to_assign_stmt_894/type_cast_880_Sample/rr
      -- CP-element group 218: 	 branch_block_stmt_26/assign_stmt_865_to_assign_stmt_894/type_cast_880_Update/$entry
      -- CP-element group 218: 	 branch_block_stmt_26/assign_stmt_865_to_assign_stmt_894/type_cast_880_Update/cr
      -- CP-element group 218: 	 branch_block_stmt_26/forx_xend250_bbx_xnph450_PhiReq/$entry
      -- CP-element group 218: 	 branch_block_stmt_26/forx_xend250_bbx_xnph450_PhiReq/$exit
      -- CP-element group 218: 	 branch_block_stmt_26/merge_stmt_859_PhiReqMerge
      -- CP-element group 218: 	 branch_block_stmt_26/merge_stmt_859_PhiAck/$entry
      -- CP-element group 218: 	 branch_block_stmt_26/merge_stmt_859_PhiAck/$exit
      -- CP-element group 218: 	 branch_block_stmt_26/merge_stmt_859_PhiAck/dummy
      -- 
    if_choice_transition_1716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_853_branch_ack_1, ack => convTranspose_CP_39_elements(218)); -- 
    rr_1733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(218), ack => type_cast_880_inst_req_0); -- 
    cr_1738_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1738_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(218), ack => type_cast_880_inst_req_1); -- 
    -- CP-element group 219:  transition  place  input  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	217 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	380 
    -- CP-element group 219:  members (5) 
      -- CP-element group 219: 	 branch_block_stmt_26/if_stmt_853_else_link/$exit
      -- CP-element group 219: 	 branch_block_stmt_26/if_stmt_853_else_link/else_choice_transition
      -- CP-element group 219: 	 branch_block_stmt_26/forx_xend250_forx_xend273
      -- CP-element group 219: 	 branch_block_stmt_26/forx_xend250_forx_xend273_PhiReq/$entry
      -- CP-element group 219: 	 branch_block_stmt_26/forx_xend250_forx_xend273_PhiReq/$exit
      -- 
    else_choice_transition_1720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_853_branch_ack_0, ack => convTranspose_CP_39_elements(219)); -- 
    -- CP-element group 220:  transition  input  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	218 
    -- CP-element group 220: successors 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_26/assign_stmt_865_to_assign_stmt_894/type_cast_880_sample_completed_
      -- CP-element group 220: 	 branch_block_stmt_26/assign_stmt_865_to_assign_stmt_894/type_cast_880_Sample/$exit
      -- CP-element group 220: 	 branch_block_stmt_26/assign_stmt_865_to_assign_stmt_894/type_cast_880_Sample/ra
      -- 
    ra_1734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_880_inst_ack_0, ack => convTranspose_CP_39_elements(220)); -- 
    -- CP-element group 221:  transition  place  input  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	218 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	374 
    -- CP-element group 221:  members (9) 
      -- CP-element group 221: 	 branch_block_stmt_26/assign_stmt_865_to_assign_stmt_894__exit__
      -- CP-element group 221: 	 branch_block_stmt_26/bbx_xnph450_forx_xbody266
      -- CP-element group 221: 	 branch_block_stmt_26/assign_stmt_865_to_assign_stmt_894/$exit
      -- CP-element group 221: 	 branch_block_stmt_26/assign_stmt_865_to_assign_stmt_894/type_cast_880_update_completed_
      -- CP-element group 221: 	 branch_block_stmt_26/assign_stmt_865_to_assign_stmt_894/type_cast_880_Update/$exit
      -- CP-element group 221: 	 branch_block_stmt_26/assign_stmt_865_to_assign_stmt_894/type_cast_880_Update/ca
      -- CP-element group 221: 	 branch_block_stmt_26/bbx_xnph450_forx_xbody266_PhiReq/$entry
      -- CP-element group 221: 	 branch_block_stmt_26/bbx_xnph450_forx_xbody266_PhiReq/phi_stmt_897/$entry
      -- CP-element group 221: 	 branch_block_stmt_26/bbx_xnph450_forx_xbody266_PhiReq/phi_stmt_897/phi_stmt_897_sources/$entry
      -- 
    ca_1739_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_880_inst_ack_1, ack => convTranspose_CP_39_elements(221)); -- 
    -- CP-element group 222:  transition  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	379 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	228 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/array_obj_ref_909_final_index_sum_regn_sample_complete
      -- CP-element group 222: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/array_obj_ref_909_final_index_sum_regn_Sample/$exit
      -- CP-element group 222: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/array_obj_ref_909_final_index_sum_regn_Sample/ack
      -- 
    ack_1768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_909_index_offset_ack_0, ack => convTranspose_CP_39_elements(222)); -- 
    -- CP-element group 223:  transition  input  output  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	379 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223:  members (11) 
      -- CP-element group 223: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/addr_of_910_sample_start_
      -- CP-element group 223: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/array_obj_ref_909_root_address_calculated
      -- CP-element group 223: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/array_obj_ref_909_offset_calculated
      -- CP-element group 223: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/array_obj_ref_909_final_index_sum_regn_Update/$exit
      -- CP-element group 223: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/array_obj_ref_909_final_index_sum_regn_Update/ack
      -- CP-element group 223: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/array_obj_ref_909_base_plus_offset/$entry
      -- CP-element group 223: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/array_obj_ref_909_base_plus_offset/$exit
      -- CP-element group 223: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/array_obj_ref_909_base_plus_offset/sum_rename_req
      -- CP-element group 223: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/array_obj_ref_909_base_plus_offset/sum_rename_ack
      -- CP-element group 223: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/addr_of_910_request/$entry
      -- CP-element group 223: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/addr_of_910_request/req
      -- 
    ack_1773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_909_index_offset_ack_1, ack => convTranspose_CP_39_elements(223)); -- 
    req_1782_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1782_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(223), ack => addr_of_910_final_reg_req_0); -- 
    -- CP-element group 224:  transition  input  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/addr_of_910_sample_completed_
      -- CP-element group 224: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/addr_of_910_request/$exit
      -- CP-element group 224: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/addr_of_910_request/ack
      -- 
    ack_1783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_910_final_reg_ack_0, ack => convTranspose_CP_39_elements(224)); -- 
    -- CP-element group 225:  join  fork  transition  input  output  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	379 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	226 
    -- CP-element group 225:  members (28) 
      -- CP-element group 225: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/addr_of_910_update_completed_
      -- CP-element group 225: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/addr_of_910_complete/$exit
      -- CP-element group 225: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/addr_of_910_complete/ack
      -- CP-element group 225: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/ptr_deref_913_sample_start_
      -- CP-element group 225: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/ptr_deref_913_base_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/ptr_deref_913_word_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/ptr_deref_913_root_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/ptr_deref_913_base_address_resized
      -- CP-element group 225: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/ptr_deref_913_base_addr_resize/$entry
      -- CP-element group 225: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/ptr_deref_913_base_addr_resize/$exit
      -- CP-element group 225: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/ptr_deref_913_base_addr_resize/base_resize_req
      -- CP-element group 225: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/ptr_deref_913_base_addr_resize/base_resize_ack
      -- CP-element group 225: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/ptr_deref_913_base_plus_offset/$entry
      -- CP-element group 225: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/ptr_deref_913_base_plus_offset/$exit
      -- CP-element group 225: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/ptr_deref_913_base_plus_offset/sum_rename_req
      -- CP-element group 225: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/ptr_deref_913_base_plus_offset/sum_rename_ack
      -- CP-element group 225: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/ptr_deref_913_word_addrgen/$entry
      -- CP-element group 225: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/ptr_deref_913_word_addrgen/$exit
      -- CP-element group 225: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/ptr_deref_913_word_addrgen/root_register_req
      -- CP-element group 225: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/ptr_deref_913_word_addrgen/root_register_ack
      -- CP-element group 225: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/ptr_deref_913_Sample/$entry
      -- CP-element group 225: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/ptr_deref_913_Sample/ptr_deref_913_Split/$entry
      -- CP-element group 225: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/ptr_deref_913_Sample/ptr_deref_913_Split/$exit
      -- CP-element group 225: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/ptr_deref_913_Sample/ptr_deref_913_Split/split_req
      -- CP-element group 225: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/ptr_deref_913_Sample/ptr_deref_913_Split/split_ack
      -- CP-element group 225: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/ptr_deref_913_Sample/word_access_start/$entry
      -- CP-element group 225: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/ptr_deref_913_Sample/word_access_start/word_0/$entry
      -- CP-element group 225: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/ptr_deref_913_Sample/word_access_start/word_0/rr
      -- 
    ack_1788_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_910_final_reg_ack_1, ack => convTranspose_CP_39_elements(225)); -- 
    rr_1826_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1826_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(225), ack => ptr_deref_913_store_0_req_0); -- 
    -- CP-element group 226:  transition  input  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	225 
    -- CP-element group 226: successors 
    -- CP-element group 226:  members (5) 
      -- CP-element group 226: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/ptr_deref_913_sample_completed_
      -- CP-element group 226: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/ptr_deref_913_Sample/$exit
      -- CP-element group 226: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/ptr_deref_913_Sample/word_access_start/$exit
      -- CP-element group 226: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/ptr_deref_913_Sample/word_access_start/word_0/$exit
      -- CP-element group 226: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/ptr_deref_913_Sample/word_access_start/word_0/ra
      -- 
    ra_1827_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_913_store_0_ack_0, ack => convTranspose_CP_39_elements(226)); -- 
    -- CP-element group 227:  transition  input  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	379 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	228 
    -- CP-element group 227:  members (5) 
      -- CP-element group 227: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/ptr_deref_913_update_completed_
      -- CP-element group 227: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/ptr_deref_913_Update/$exit
      -- CP-element group 227: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/ptr_deref_913_Update/word_access_complete/$exit
      -- CP-element group 227: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/ptr_deref_913_Update/word_access_complete/word_0/$exit
      -- CP-element group 227: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/ptr_deref_913_Update/word_access_complete/word_0/ca
      -- 
    ca_1838_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_913_store_0_ack_1, ack => convTranspose_CP_39_elements(227)); -- 
    -- CP-element group 228:  branch  join  transition  place  output  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	222 
    -- CP-element group 228: 	227 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	229 
    -- CP-element group 228: 	230 
    -- CP-element group 228:  members (10) 
      -- CP-element group 228: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927__exit__
      -- CP-element group 228: 	 branch_block_stmt_26/if_stmt_928__entry__
      -- CP-element group 228: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/$exit
      -- CP-element group 228: 	 branch_block_stmt_26/if_stmt_928_dead_link/$entry
      -- CP-element group 228: 	 branch_block_stmt_26/if_stmt_928_eval_test/$entry
      -- CP-element group 228: 	 branch_block_stmt_26/if_stmt_928_eval_test/$exit
      -- CP-element group 228: 	 branch_block_stmt_26/if_stmt_928_eval_test/branch_req
      -- CP-element group 228: 	 branch_block_stmt_26/R_exitcond_929_place
      -- CP-element group 228: 	 branch_block_stmt_26/if_stmt_928_if_link/$entry
      -- CP-element group 228: 	 branch_block_stmt_26/if_stmt_928_else_link/$entry
      -- 
    branch_req_1846_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1846_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(228), ack => if_stmt_928_branch_req_0); -- 
    convTranspose_cp_element_group_228: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_228"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(222) & convTranspose_CP_39_elements(227);
      gj_convTranspose_cp_element_group_228 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(228), clk => clk, reset => reset); --
    end block;
    -- CP-element group 229:  merge  transition  place  input  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	228 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	380 
    -- CP-element group 229:  members (13) 
      -- CP-element group 229: 	 branch_block_stmt_26/merge_stmt_934__exit__
      -- CP-element group 229: 	 branch_block_stmt_26/forx_xend273x_xloopexit_forx_xend273
      -- CP-element group 229: 	 branch_block_stmt_26/if_stmt_928_if_link/$exit
      -- CP-element group 229: 	 branch_block_stmt_26/if_stmt_928_if_link/if_choice_transition
      -- CP-element group 229: 	 branch_block_stmt_26/forx_xbody266_forx_xend273x_xloopexit
      -- CP-element group 229: 	 branch_block_stmt_26/forx_xbody266_forx_xend273x_xloopexit_PhiReq/$entry
      -- CP-element group 229: 	 branch_block_stmt_26/forx_xbody266_forx_xend273x_xloopexit_PhiReq/$exit
      -- CP-element group 229: 	 branch_block_stmt_26/merge_stmt_934_PhiReqMerge
      -- CP-element group 229: 	 branch_block_stmt_26/merge_stmt_934_PhiAck/$entry
      -- CP-element group 229: 	 branch_block_stmt_26/merge_stmt_934_PhiAck/$exit
      -- CP-element group 229: 	 branch_block_stmt_26/merge_stmt_934_PhiAck/dummy
      -- CP-element group 229: 	 branch_block_stmt_26/forx_xend273x_xloopexit_forx_xend273_PhiReq/$entry
      -- CP-element group 229: 	 branch_block_stmt_26/forx_xend273x_xloopexit_forx_xend273_PhiReq/$exit
      -- 
    if_choice_transition_1851_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_928_branch_ack_1, ack => convTranspose_CP_39_elements(229)); -- 
    -- CP-element group 230:  fork  transition  place  input  output  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	228 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	375 
    -- CP-element group 230: 	376 
    -- CP-element group 230:  members (12) 
      -- CP-element group 230: 	 branch_block_stmt_26/if_stmt_928_else_link/$exit
      -- CP-element group 230: 	 branch_block_stmt_26/if_stmt_928_else_link/else_choice_transition
      -- CP-element group 230: 	 branch_block_stmt_26/forx_xbody266_forx_xbody266
      -- CP-element group 230: 	 branch_block_stmt_26/forx_xbody266_forx_xbody266_PhiReq/$entry
      -- CP-element group 230: 	 branch_block_stmt_26/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_897/$entry
      -- CP-element group 230: 	 branch_block_stmt_26/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_897/phi_stmt_897_sources/$entry
      -- CP-element group 230: 	 branch_block_stmt_26/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_897/phi_stmt_897_sources/type_cast_903/$entry
      -- CP-element group 230: 	 branch_block_stmt_26/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_897/phi_stmt_897_sources/type_cast_903/SplitProtocol/$entry
      -- CP-element group 230: 	 branch_block_stmt_26/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_897/phi_stmt_897_sources/type_cast_903/SplitProtocol/Sample/$entry
      -- CP-element group 230: 	 branch_block_stmt_26/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_897/phi_stmt_897_sources/type_cast_903/SplitProtocol/Sample/rr
      -- CP-element group 230: 	 branch_block_stmt_26/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_897/phi_stmt_897_sources/type_cast_903/SplitProtocol/Update/$entry
      -- CP-element group 230: 	 branch_block_stmt_26/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_897/phi_stmt_897_sources/type_cast_903/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_928_branch_ack_0, ack => convTranspose_CP_39_elements(230)); -- 
    rr_2933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(230), ack => type_cast_903_inst_req_0); -- 
    cr_2938_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2938_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(230), ack => type_cast_903_inst_req_1); -- 
    -- CP-element group 231:  transition  input  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	380 
    -- CP-element group 231: successors 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 branch_block_stmt_26/call_stmt_939_to_assign_stmt_945/call_stmt_939_sample_completed_
      -- CP-element group 231: 	 branch_block_stmt_26/call_stmt_939_to_assign_stmt_945/call_stmt_939_Sample/$exit
      -- CP-element group 231: 	 branch_block_stmt_26/call_stmt_939_to_assign_stmt_945/call_stmt_939_Sample/cra
      -- 
    cra_1869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_939_call_ack_0, ack => convTranspose_CP_39_elements(231)); -- 
    -- CP-element group 232:  transition  input  output  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	380 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	233 
    -- CP-element group 232:  members (6) 
      -- CP-element group 232: 	 branch_block_stmt_26/call_stmt_939_to_assign_stmt_945/call_stmt_939_update_completed_
      -- CP-element group 232: 	 branch_block_stmt_26/call_stmt_939_to_assign_stmt_945/call_stmt_939_Update/$exit
      -- CP-element group 232: 	 branch_block_stmt_26/call_stmt_939_to_assign_stmt_945/call_stmt_939_Update/cca
      -- CP-element group 232: 	 branch_block_stmt_26/call_stmt_939_to_assign_stmt_945/type_cast_944_sample_start_
      -- CP-element group 232: 	 branch_block_stmt_26/call_stmt_939_to_assign_stmt_945/type_cast_944_Sample/$entry
      -- CP-element group 232: 	 branch_block_stmt_26/call_stmt_939_to_assign_stmt_945/type_cast_944_Sample/rr
      -- 
    cca_1874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_939_call_ack_1, ack => convTranspose_CP_39_elements(232)); -- 
    rr_1882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(232), ack => type_cast_944_inst_req_0); -- 
    -- CP-element group 233:  transition  input  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	232 
    -- CP-element group 233: successors 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_26/call_stmt_939_to_assign_stmt_945/type_cast_944_sample_completed_
      -- CP-element group 233: 	 branch_block_stmt_26/call_stmt_939_to_assign_stmt_945/type_cast_944_Sample/$exit
      -- CP-element group 233: 	 branch_block_stmt_26/call_stmt_939_to_assign_stmt_945/type_cast_944_Sample/ra
      -- 
    ra_1883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_944_inst_ack_0, ack => convTranspose_CP_39_elements(233)); -- 
    -- CP-element group 234:  transition  place  input  output  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	380 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	235 
    -- CP-element group 234:  members (10) 
      -- CP-element group 234: 	 branch_block_stmt_26/call_stmt_939_to_assign_stmt_945__exit__
      -- CP-element group 234: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990__entry__
      -- CP-element group 234: 	 branch_block_stmt_26/call_stmt_939_to_assign_stmt_945/$exit
      -- CP-element group 234: 	 branch_block_stmt_26/call_stmt_939_to_assign_stmt_945/type_cast_944_update_completed_
      -- CP-element group 234: 	 branch_block_stmt_26/call_stmt_939_to_assign_stmt_945/type_cast_944_Update/$exit
      -- CP-element group 234: 	 branch_block_stmt_26/call_stmt_939_to_assign_stmt_945/type_cast_944_Update/ca
      -- CP-element group 234: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/$entry
      -- CP-element group 234: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_947_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_947_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_947_Sample/req
      -- 
    ca_1888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_944_inst_ack_1, ack => convTranspose_CP_39_elements(234)); -- 
    req_1899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => WPIPE_Block0_start_947_inst_req_0); -- 
    -- CP-element group 235:  transition  input  output  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	234 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235:  members (6) 
      -- CP-element group 235: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_947_sample_completed_
      -- CP-element group 235: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_947_update_start_
      -- CP-element group 235: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_947_Sample/$exit
      -- CP-element group 235: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_947_Sample/ack
      -- CP-element group 235: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_947_Update/$entry
      -- CP-element group 235: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_947_Update/req
      -- 
    ack_1900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_947_inst_ack_0, ack => convTranspose_CP_39_elements(235)); -- 
    req_1904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(235), ack => WPIPE_Block0_start_947_inst_req_1); -- 
    -- CP-element group 236:  transition  input  output  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	237 
    -- CP-element group 236:  members (6) 
      -- CP-element group 236: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_947_update_completed_
      -- CP-element group 236: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_947_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_947_Update/ack
      -- CP-element group 236: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_950_sample_start_
      -- CP-element group 236: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_950_Sample/$entry
      -- CP-element group 236: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_950_Sample/req
      -- 
    ack_1905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_947_inst_ack_1, ack => convTranspose_CP_39_elements(236)); -- 
    req_1913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(236), ack => WPIPE_Block0_start_950_inst_req_0); -- 
    -- CP-element group 237:  transition  input  output  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	236 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	238 
    -- CP-element group 237:  members (6) 
      -- CP-element group 237: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_950_Update/req
      -- CP-element group 237: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_950_Update/$entry
      -- CP-element group 237: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_950_Sample/ack
      -- CP-element group 237: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_950_sample_completed_
      -- CP-element group 237: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_950_update_start_
      -- CP-element group 237: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_950_Sample/$exit
      -- 
    ack_1914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_950_inst_ack_0, ack => convTranspose_CP_39_elements(237)); -- 
    req_1918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(237), ack => WPIPE_Block0_start_950_inst_req_1); -- 
    -- CP-element group 238:  transition  input  output  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	237 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	239 
    -- CP-element group 238:  members (6) 
      -- CP-element group 238: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_950_Update/$exit
      -- CP-element group 238: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_950_Update/ack
      -- CP-element group 238: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_953_sample_start_
      -- CP-element group 238: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_953_Sample/req
      -- CP-element group 238: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_953_Sample/$entry
      -- CP-element group 238: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_950_update_completed_
      -- 
    ack_1919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_950_inst_ack_1, ack => convTranspose_CP_39_elements(238)); -- 
    req_1927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(238), ack => WPIPE_Block0_start_953_inst_req_0); -- 
    -- CP-element group 239:  transition  input  output  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	238 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	240 
    -- CP-element group 239:  members (6) 
      -- CP-element group 239: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_953_Update/req
      -- CP-element group 239: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_953_update_start_
      -- CP-element group 239: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_953_Update/$entry
      -- CP-element group 239: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_953_Sample/$exit
      -- CP-element group 239: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_953_Sample/ack
      -- CP-element group 239: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_953_sample_completed_
      -- 
    ack_1928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_953_inst_ack_0, ack => convTranspose_CP_39_elements(239)); -- 
    req_1932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(239), ack => WPIPE_Block0_start_953_inst_req_1); -- 
    -- CP-element group 240:  transition  input  output  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	239 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	241 
    -- CP-element group 240:  members (6) 
      -- CP-element group 240: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_953_Update/$exit
      -- CP-element group 240: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_953_update_completed_
      -- CP-element group 240: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_953_Update/ack
      -- CP-element group 240: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_956_sample_start_
      -- CP-element group 240: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_956_Sample/$entry
      -- CP-element group 240: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_956_Sample/req
      -- 
    ack_1933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_953_inst_ack_1, ack => convTranspose_CP_39_elements(240)); -- 
    req_1941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(240), ack => WPIPE_Block0_start_956_inst_req_0); -- 
    -- CP-element group 241:  transition  input  output  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	240 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	242 
    -- CP-element group 241:  members (6) 
      -- CP-element group 241: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_956_sample_completed_
      -- CP-element group 241: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_956_update_start_
      -- CP-element group 241: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_956_Sample/$exit
      -- CP-element group 241: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_956_Update/req
      -- CP-element group 241: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_956_Update/$entry
      -- CP-element group 241: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_956_Sample/ack
      -- 
    ack_1942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_956_inst_ack_0, ack => convTranspose_CP_39_elements(241)); -- 
    req_1946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(241), ack => WPIPE_Block0_start_956_inst_req_1); -- 
    -- CP-element group 242:  transition  input  output  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	241 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	243 
    -- CP-element group 242:  members (6) 
      -- CP-element group 242: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_956_update_completed_
      -- CP-element group 242: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_959_Sample/req
      -- CP-element group 242: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_959_Sample/$entry
      -- CP-element group 242: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_959_sample_start_
      -- CP-element group 242: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_956_Update/ack
      -- CP-element group 242: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_956_Update/$exit
      -- 
    ack_1947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_956_inst_ack_1, ack => convTranspose_CP_39_elements(242)); -- 
    req_1955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(242), ack => WPIPE_Block0_start_959_inst_req_0); -- 
    -- CP-element group 243:  transition  input  output  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	242 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	244 
    -- CP-element group 243:  members (6) 
      -- CP-element group 243: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_959_Update/$entry
      -- CP-element group 243: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_959_Update/req
      -- CP-element group 243: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_959_Sample/ack
      -- CP-element group 243: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_959_Sample/$exit
      -- CP-element group 243: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_959_update_start_
      -- CP-element group 243: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_959_sample_completed_
      -- 
    ack_1956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_959_inst_ack_0, ack => convTranspose_CP_39_elements(243)); -- 
    req_1960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(243), ack => WPIPE_Block0_start_959_inst_req_1); -- 
    -- CP-element group 244:  transition  input  output  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	243 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	245 
    -- CP-element group 244:  members (6) 
      -- CP-element group 244: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_959_Update/$exit
      -- CP-element group 244: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_962_Sample/req
      -- CP-element group 244: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_962_sample_start_
      -- CP-element group 244: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_959_Update/ack
      -- CP-element group 244: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_962_Sample/$entry
      -- CP-element group 244: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_959_update_completed_
      -- 
    ack_1961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_959_inst_ack_1, ack => convTranspose_CP_39_elements(244)); -- 
    req_1969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(244), ack => WPIPE_Block0_start_962_inst_req_0); -- 
    -- CP-element group 245:  transition  input  output  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	244 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	246 
    -- CP-element group 245:  members (6) 
      -- CP-element group 245: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_962_update_start_
      -- CP-element group 245: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_962_sample_completed_
      -- CP-element group 245: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_962_Sample/$exit
      -- CP-element group 245: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_962_Update/req
      -- CP-element group 245: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_962_Update/$entry
      -- CP-element group 245: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_962_Sample/ack
      -- 
    ack_1970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_962_inst_ack_0, ack => convTranspose_CP_39_elements(245)); -- 
    req_1974_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1974_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(245), ack => WPIPE_Block0_start_962_inst_req_1); -- 
    -- CP-element group 246:  transition  input  output  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	245 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	247 
    -- CP-element group 246:  members (6) 
      -- CP-element group 246: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_962_update_completed_
      -- CP-element group 246: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_965_Sample/req
      -- CP-element group 246: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_965_Sample/$entry
      -- CP-element group 246: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_965_sample_start_
      -- CP-element group 246: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_962_Update/ack
      -- CP-element group 246: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_962_Update/$exit
      -- 
    ack_1975_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_962_inst_ack_1, ack => convTranspose_CP_39_elements(246)); -- 
    req_1983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(246), ack => WPIPE_Block0_start_965_inst_req_0); -- 
    -- CP-element group 247:  transition  input  output  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	246 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	248 
    -- CP-element group 247:  members (6) 
      -- CP-element group 247: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_965_Update/req
      -- CP-element group 247: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_965_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_965_Sample/ack
      -- CP-element group 247: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_965_Sample/$exit
      -- CP-element group 247: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_965_update_start_
      -- CP-element group 247: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_965_sample_completed_
      -- 
    ack_1984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_965_inst_ack_0, ack => convTranspose_CP_39_elements(247)); -- 
    req_1988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(247), ack => WPIPE_Block0_start_965_inst_req_1); -- 
    -- CP-element group 248:  transition  input  output  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	247 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	249 
    -- CP-element group 248:  members (6) 
      -- CP-element group 248: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_965_Update/$exit
      -- CP-element group 248: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_968_Sample/req
      -- CP-element group 248: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_965_Update/ack
      -- CP-element group 248: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_968_sample_start_
      -- CP-element group 248: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_968_Sample/$entry
      -- CP-element group 248: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_965_update_completed_
      -- 
    ack_1989_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_965_inst_ack_1, ack => convTranspose_CP_39_elements(248)); -- 
    req_1997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(248), ack => WPIPE_Block0_start_968_inst_req_0); -- 
    -- CP-element group 249:  transition  input  output  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	248 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	250 
    -- CP-element group 249:  members (6) 
      -- CP-element group 249: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_968_Sample/$exit
      -- CP-element group 249: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_968_update_start_
      -- CP-element group 249: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_968_sample_completed_
      -- CP-element group 249: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_968_Update/req
      -- CP-element group 249: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_968_Sample/ack
      -- CP-element group 249: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_968_Update/$entry
      -- 
    ack_1998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_968_inst_ack_0, ack => convTranspose_CP_39_elements(249)); -- 
    req_2002_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2002_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(249), ack => WPIPE_Block0_start_968_inst_req_1); -- 
    -- CP-element group 250:  transition  input  output  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	249 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	251 
    -- CP-element group 250:  members (6) 
      -- CP-element group 250: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_968_Update/$exit
      -- CP-element group 250: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_968_update_completed_
      -- CP-element group 250: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_968_Update/ack
      -- CP-element group 250: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_971_sample_start_
      -- CP-element group 250: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_971_Sample/$entry
      -- CP-element group 250: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_971_Sample/req
      -- 
    ack_2003_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_968_inst_ack_1, ack => convTranspose_CP_39_elements(250)); -- 
    req_2011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(250), ack => WPIPE_Block0_start_971_inst_req_0); -- 
    -- CP-element group 251:  transition  input  output  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	250 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	252 
    -- CP-element group 251:  members (6) 
      -- CP-element group 251: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_971_sample_completed_
      -- CP-element group 251: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_971_update_start_
      -- CP-element group 251: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_971_Sample/$exit
      -- CP-element group 251: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_971_Sample/ack
      -- CP-element group 251: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_971_Update/$entry
      -- CP-element group 251: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_971_Update/req
      -- 
    ack_2012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_971_inst_ack_0, ack => convTranspose_CP_39_elements(251)); -- 
    req_2016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(251), ack => WPIPE_Block0_start_971_inst_req_1); -- 
    -- CP-element group 252:  transition  input  output  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	251 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	253 
    -- CP-element group 252:  members (6) 
      -- CP-element group 252: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_971_update_completed_
      -- CP-element group 252: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_971_Update/$exit
      -- CP-element group 252: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_971_Update/ack
      -- CP-element group 252: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_974_sample_start_
      -- CP-element group 252: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_974_Sample/req
      -- CP-element group 252: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_974_Sample/$entry
      -- 
    ack_2017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_971_inst_ack_1, ack => convTranspose_CP_39_elements(252)); -- 
    req_2025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(252), ack => WPIPE_Block0_start_974_inst_req_0); -- 
    -- CP-element group 253:  transition  input  output  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	252 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	254 
    -- CP-element group 253:  members (6) 
      -- CP-element group 253: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_974_sample_completed_
      -- CP-element group 253: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_974_update_start_
      -- CP-element group 253: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_974_Update/req
      -- CP-element group 253: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_974_Update/$entry
      -- CP-element group 253: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_974_Sample/ack
      -- CP-element group 253: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_974_Sample/$exit
      -- 
    ack_2026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_974_inst_ack_0, ack => convTranspose_CP_39_elements(253)); -- 
    req_2030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(253), ack => WPIPE_Block0_start_974_inst_req_1); -- 
    -- CP-element group 254:  transition  input  output  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	253 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	255 
    -- CP-element group 254:  members (6) 
      -- CP-element group 254: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_978_sample_start_
      -- CP-element group 254: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_978_Sample/$entry
      -- CP-element group 254: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_978_Sample/req
      -- CP-element group 254: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_974_Update/ack
      -- CP-element group 254: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_974_Update/$exit
      -- CP-element group 254: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_974_update_completed_
      -- 
    ack_2031_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_974_inst_ack_1, ack => convTranspose_CP_39_elements(254)); -- 
    req_2039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(254), ack => WPIPE_Block0_start_978_inst_req_0); -- 
    -- CP-element group 255:  transition  input  output  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	254 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	256 
    -- CP-element group 255:  members (6) 
      -- CP-element group 255: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_978_update_start_
      -- CP-element group 255: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_978_sample_completed_
      -- CP-element group 255: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_978_Update/$entry
      -- CP-element group 255: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_978_Sample/$exit
      -- CP-element group 255: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_978_Sample/ack
      -- CP-element group 255: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_978_Update/req
      -- 
    ack_2040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_978_inst_ack_0, ack => convTranspose_CP_39_elements(255)); -- 
    req_2044_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2044_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(255), ack => WPIPE_Block0_start_978_inst_req_1); -- 
    -- CP-element group 256:  transition  input  output  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	255 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	257 
    -- CP-element group 256:  members (6) 
      -- CP-element group 256: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_978_update_completed_
      -- CP-element group 256: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_982_Sample/req
      -- CP-element group 256: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_982_Sample/$entry
      -- CP-element group 256: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_982_sample_start_
      -- CP-element group 256: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_978_Update/ack
      -- CP-element group 256: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_978_Update/$exit
      -- 
    ack_2045_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_978_inst_ack_1, ack => convTranspose_CP_39_elements(256)); -- 
    req_2053_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2053_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(256), ack => WPIPE_Block0_start_982_inst_req_0); -- 
    -- CP-element group 257:  transition  input  output  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	256 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	258 
    -- CP-element group 257:  members (6) 
      -- CP-element group 257: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_982_Update/req
      -- CP-element group 257: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_982_Update/$entry
      -- CP-element group 257: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_982_Sample/ack
      -- CP-element group 257: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_982_Sample/$exit
      -- CP-element group 257: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_982_update_start_
      -- CP-element group 257: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_982_sample_completed_
      -- 
    ack_2054_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_982_inst_ack_0, ack => convTranspose_CP_39_elements(257)); -- 
    req_2058_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2058_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(257), ack => WPIPE_Block0_start_982_inst_req_1); -- 
    -- CP-element group 258:  transition  input  output  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	257 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	259 
    -- CP-element group 258:  members (6) 
      -- CP-element group 258: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_985_Sample/req
      -- CP-element group 258: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_985_Sample/$entry
      -- CP-element group 258: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_985_sample_start_
      -- CP-element group 258: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_982_Update/ack
      -- CP-element group 258: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_982_Update/$exit
      -- CP-element group 258: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_982_update_completed_
      -- 
    ack_2059_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_982_inst_ack_1, ack => convTranspose_CP_39_elements(258)); -- 
    req_2067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(258), ack => WPIPE_Block0_start_985_inst_req_0); -- 
    -- CP-element group 259:  transition  input  output  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	258 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	260 
    -- CP-element group 259:  members (6) 
      -- CP-element group 259: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_985_Update/req
      -- CP-element group 259: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_985_Update/$entry
      -- CP-element group 259: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_985_Sample/ack
      -- CP-element group 259: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_985_Sample/$exit
      -- CP-element group 259: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_985_update_start_
      -- CP-element group 259: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_985_sample_completed_
      -- 
    ack_2068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_985_inst_ack_0, ack => convTranspose_CP_39_elements(259)); -- 
    req_2072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(259), ack => WPIPE_Block0_start_985_inst_req_1); -- 
    -- CP-element group 260:  transition  input  output  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	259 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	261 
    -- CP-element group 260:  members (6) 
      -- CP-element group 260: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_988_Sample/req
      -- CP-element group 260: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_988_Sample/$entry
      -- CP-element group 260: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_988_sample_start_
      -- CP-element group 260: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_985_Update/ack
      -- CP-element group 260: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_985_Update/$exit
      -- CP-element group 260: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_985_update_completed_
      -- 
    ack_2073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_985_inst_ack_1, ack => convTranspose_CP_39_elements(260)); -- 
    req_2081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(260), ack => WPIPE_Block0_start_988_inst_req_0); -- 
    -- CP-element group 261:  transition  input  output  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	260 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	262 
    -- CP-element group 261:  members (6) 
      -- CP-element group 261: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_988_Update/$entry
      -- CP-element group 261: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_988_Update/req
      -- CP-element group 261: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_988_Sample/ack
      -- CP-element group 261: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_988_Sample/$exit
      -- CP-element group 261: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_988_update_start_
      -- CP-element group 261: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_988_sample_completed_
      -- 
    ack_2082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_988_inst_ack_0, ack => convTranspose_CP_39_elements(261)); -- 
    req_2086_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2086_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(261), ack => WPIPE_Block0_start_988_inst_req_1); -- 
    -- CP-element group 262:  transition  place  input  output  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	261 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	263 
    -- CP-element group 262:  members (10) 
      -- CP-element group 262: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_988_Update/$exit
      -- CP-element group 262: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990__exit__
      -- CP-element group 262: 	 branch_block_stmt_26/assign_stmt_994__entry__
      -- CP-element group 262: 	 branch_block_stmt_26/assign_stmt_994/RPIPE_Block0_done_993_Sample/$entry
      -- CP-element group 262: 	 branch_block_stmt_26/assign_stmt_994/RPIPE_Block0_done_993_Sample/rr
      -- CP-element group 262: 	 branch_block_stmt_26/assign_stmt_994/RPIPE_Block0_done_993_sample_start_
      -- CP-element group 262: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_988_Update/ack
      -- CP-element group 262: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/WPIPE_Block0_start_988_update_completed_
      -- CP-element group 262: 	 branch_block_stmt_26/assign_stmt_994/$entry
      -- CP-element group 262: 	 branch_block_stmt_26/assign_stmt_949_to_assign_stmt_990/$exit
      -- 
    ack_2087_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_988_inst_ack_1, ack => convTranspose_CP_39_elements(262)); -- 
    rr_2098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(262), ack => RPIPE_Block0_done_993_inst_req_0); -- 
    -- CP-element group 263:  transition  input  output  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	262 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	264 
    -- CP-element group 263:  members (6) 
      -- CP-element group 263: 	 branch_block_stmt_26/assign_stmt_994/RPIPE_Block0_done_993_sample_completed_
      -- CP-element group 263: 	 branch_block_stmt_26/assign_stmt_994/RPIPE_Block0_done_993_Sample/ra
      -- CP-element group 263: 	 branch_block_stmt_26/assign_stmt_994/RPIPE_Block0_done_993_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_26/assign_stmt_994/RPIPE_Block0_done_993_Sample/$exit
      -- CP-element group 263: 	 branch_block_stmt_26/assign_stmt_994/RPIPE_Block0_done_993_Update/cr
      -- CP-element group 263: 	 branch_block_stmt_26/assign_stmt_994/RPIPE_Block0_done_993_update_start_
      -- 
    ra_2099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_993_inst_ack_0, ack => convTranspose_CP_39_elements(263)); -- 
    cr_2103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(263), ack => RPIPE_Block0_done_993_inst_req_1); -- 
    -- CP-element group 264:  fork  transition  place  input  output  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	263 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	265 
    -- CP-element group 264: 	266 
    -- CP-element group 264: 	268 
    -- CP-element group 264: 	270 
    -- CP-element group 264: 	272 
    -- CP-element group 264: 	274 
    -- CP-element group 264: 	276 
    -- CP-element group 264: 	278 
    -- CP-element group 264: 	280 
    -- CP-element group 264: 	282 
    -- CP-element group 264: 	284 
    -- CP-element group 264:  members (40) 
      -- CP-element group 264: 	 branch_block_stmt_26/assign_stmt_994/RPIPE_Block0_done_993_update_completed_
      -- CP-element group 264: 	 branch_block_stmt_26/assign_stmt_994__exit__
      -- CP-element group 264: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105__entry__
      -- CP-element group 264: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1060_Update/$entry
      -- CP-element group 264: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1060_Update/cr
      -- CP-element group 264: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/call_stmt_997_Sample/crr
      -- CP-element group 264: 	 branch_block_stmt_26/assign_stmt_994/RPIPE_Block0_done_993_Update/$exit
      -- CP-element group 264: 	 branch_block_stmt_26/assign_stmt_994/$exit
      -- CP-element group 264: 	 branch_block_stmt_26/assign_stmt_994/RPIPE_Block0_done_993_Update/ca
      -- CP-element group 264: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1001_update_start_
      -- CP-element group 264: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/$entry
      -- CP-element group 264: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/call_stmt_997_sample_start_
      -- CP-element group 264: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/call_stmt_997_update_start_
      -- CP-element group 264: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1070_Update/$entry
      -- CP-element group 264: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1070_update_start_
      -- CP-element group 264: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/call_stmt_997_Sample/$entry
      -- CP-element group 264: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/call_stmt_997_Update/$entry
      -- CP-element group 264: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/call_stmt_997_Update/ccr
      -- CP-element group 264: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1060_update_start_
      -- CP-element group 264: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1080_Update/cr
      -- CP-element group 264: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1050_Update/cr
      -- CP-element group 264: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1080_Update/$entry
      -- CP-element group 264: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1050_Update/$entry
      -- CP-element group 264: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1050_update_start_
      -- CP-element group 264: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1020_update_start_
      -- CP-element group 264: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1040_Update/cr
      -- CP-element group 264: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1010_Update/cr
      -- CP-element group 264: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1010_Update/$entry
      -- CP-element group 264: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1080_update_start_
      -- CP-element group 264: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1040_Update/$entry
      -- CP-element group 264: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1010_update_start_
      -- CP-element group 264: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1040_update_start_
      -- CP-element group 264: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1030_Update/cr
      -- CP-element group 264: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1030_Update/$entry
      -- CP-element group 264: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1001_Update/cr
      -- CP-element group 264: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1001_Update/$entry
      -- CP-element group 264: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1030_update_start_
      -- CP-element group 264: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1070_Update/cr
      -- CP-element group 264: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1020_Update/cr
      -- CP-element group 264: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1020_Update/$entry
      -- 
    ca_2104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_993_inst_ack_1, ack => convTranspose_CP_39_elements(264)); -- 
    cr_2218_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2218_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(264), ack => type_cast_1060_inst_req_1); -- 
    crr_2115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(264), ack => call_stmt_997_call_req_0); -- 
    ccr_2120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(264), ack => call_stmt_997_call_req_1); -- 
    cr_2246_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2246_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(264), ack => type_cast_1080_inst_req_1); -- 
    cr_2204_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2204_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(264), ack => type_cast_1050_inst_req_1); -- 
    cr_2190_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2190_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(264), ack => type_cast_1040_inst_req_1); -- 
    cr_2148_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2148_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(264), ack => type_cast_1010_inst_req_1); -- 
    cr_2176_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2176_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(264), ack => type_cast_1030_inst_req_1); -- 
    cr_2134_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2134_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(264), ack => type_cast_1001_inst_req_1); -- 
    cr_2232_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2232_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(264), ack => type_cast_1070_inst_req_1); -- 
    cr_2162_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2162_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(264), ack => type_cast_1020_inst_req_1); -- 
    -- CP-element group 265:  transition  input  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	264 
    -- CP-element group 265: successors 
    -- CP-element group 265:  members (3) 
      -- CP-element group 265: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/call_stmt_997_sample_completed_
      -- CP-element group 265: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/call_stmt_997_Sample/$exit
      -- CP-element group 265: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/call_stmt_997_Sample/cra
      -- 
    cra_2116_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_997_call_ack_0, ack => convTranspose_CP_39_elements(265)); -- 
    -- CP-element group 266:  transition  input  output  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	264 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	267 
    -- CP-element group 266:  members (6) 
      -- CP-element group 266: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/call_stmt_997_update_completed_
      -- CP-element group 266: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/call_stmt_997_Update/$exit
      -- CP-element group 266: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/call_stmt_997_Update/cca
      -- CP-element group 266: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1001_sample_start_
      -- CP-element group 266: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1001_Sample/rr
      -- CP-element group 266: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1001_Sample/$entry
      -- 
    cca_2121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_997_call_ack_1, ack => convTranspose_CP_39_elements(266)); -- 
    rr_2129_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2129_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(266), ack => type_cast_1001_inst_req_0); -- 
    -- CP-element group 267:  transition  input  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	266 
    -- CP-element group 267: successors 
    -- CP-element group 267:  members (3) 
      -- CP-element group 267: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1001_sample_completed_
      -- CP-element group 267: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1001_Sample/ra
      -- CP-element group 267: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1001_Sample/$exit
      -- 
    ra_2130_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1001_inst_ack_0, ack => convTranspose_CP_39_elements(267)); -- 
    -- CP-element group 268:  fork  transition  input  output  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	264 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	269 
    -- CP-element group 268: 	271 
    -- CP-element group 268: 	273 
    -- CP-element group 268: 	275 
    -- CP-element group 268: 	277 
    -- CP-element group 268: 	279 
    -- CP-element group 268: 	281 
    -- CP-element group 268: 	283 
    -- CP-element group 268:  members (27) 
      -- CP-element group 268: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1060_Sample/rr
      -- CP-element group 268: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1020_Sample/$entry
      -- CP-element group 268: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1070_sample_start_
      -- CP-element group 268: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1020_Sample/rr
      -- CP-element group 268: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1070_Sample/$entry
      -- CP-element group 268: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1070_Sample/rr
      -- CP-element group 268: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1060_Sample/$entry
      -- CP-element group 268: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1060_sample_start_
      -- CP-element group 268: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1050_Sample/rr
      -- CP-element group 268: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1050_Sample/$entry
      -- CP-element group 268: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1080_Sample/rr
      -- CP-element group 268: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1080_Sample/$entry
      -- CP-element group 268: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1050_sample_start_
      -- CP-element group 268: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1020_sample_start_
      -- CP-element group 268: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1040_Sample/rr
      -- CP-element group 268: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1080_sample_start_
      -- CP-element group 268: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1040_Sample/$entry
      -- CP-element group 268: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1010_Sample/rr
      -- CP-element group 268: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1010_Sample/$entry
      -- CP-element group 268: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1010_sample_start_
      -- CP-element group 268: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1001_Update/ca
      -- CP-element group 268: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1040_sample_start_
      -- CP-element group 268: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1030_Sample/rr
      -- CP-element group 268: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1030_Sample/$entry
      -- CP-element group 268: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1001_Update/$exit
      -- CP-element group 268: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1030_sample_start_
      -- CP-element group 268: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1001_update_completed_
      -- 
    ca_2135_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1001_inst_ack_1, ack => convTranspose_CP_39_elements(268)); -- 
    rr_2143_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2143_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(268), ack => type_cast_1010_inst_req_0); -- 
    rr_2157_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2157_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(268), ack => type_cast_1020_inst_req_0); -- 
    rr_2171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(268), ack => type_cast_1030_inst_req_0); -- 
    rr_2185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(268), ack => type_cast_1040_inst_req_0); -- 
    rr_2199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(268), ack => type_cast_1050_inst_req_0); -- 
    rr_2213_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2213_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(268), ack => type_cast_1060_inst_req_0); -- 
    rr_2227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(268), ack => type_cast_1070_inst_req_0); -- 
    rr_2241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(268), ack => type_cast_1080_inst_req_0); -- 
    -- CP-element group 269:  transition  input  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	268 
    -- CP-element group 269: successors 
    -- CP-element group 269:  members (3) 
      -- CP-element group 269: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1010_Sample/ra
      -- CP-element group 269: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1010_Sample/$exit
      -- CP-element group 269: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1010_sample_completed_
      -- 
    ra_2144_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 269_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1010_inst_ack_0, ack => convTranspose_CP_39_elements(269)); -- 
    -- CP-element group 270:  transition  input  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	264 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	305 
    -- CP-element group 270:  members (3) 
      -- CP-element group 270: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1010_Update/ca
      -- CP-element group 270: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1010_Update/$exit
      -- CP-element group 270: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1010_update_completed_
      -- 
    ca_2149_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1010_inst_ack_1, ack => convTranspose_CP_39_elements(270)); -- 
    -- CP-element group 271:  transition  input  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	268 
    -- CP-element group 271: successors 
    -- CP-element group 271:  members (3) 
      -- CP-element group 271: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1020_Sample/$exit
      -- CP-element group 271: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1020_Sample/ra
      -- CP-element group 271: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1020_sample_completed_
      -- 
    ra_2158_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1020_inst_ack_0, ack => convTranspose_CP_39_elements(271)); -- 
    -- CP-element group 272:  transition  input  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	264 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	302 
    -- CP-element group 272:  members (3) 
      -- CP-element group 272: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1020_update_completed_
      -- CP-element group 272: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1020_Update/ca
      -- CP-element group 272: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1020_Update/$exit
      -- 
    ca_2163_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1020_inst_ack_1, ack => convTranspose_CP_39_elements(272)); -- 
    -- CP-element group 273:  transition  input  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	268 
    -- CP-element group 273: successors 
    -- CP-element group 273:  members (3) 
      -- CP-element group 273: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1030_Sample/ra
      -- CP-element group 273: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1030_Sample/$exit
      -- CP-element group 273: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1030_sample_completed_
      -- 
    ra_2172_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1030_inst_ack_0, ack => convTranspose_CP_39_elements(273)); -- 
    -- CP-element group 274:  transition  input  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	264 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	299 
    -- CP-element group 274:  members (3) 
      -- CP-element group 274: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1030_Update/ca
      -- CP-element group 274: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1030_Update/$exit
      -- CP-element group 274: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1030_update_completed_
      -- 
    ca_2177_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1030_inst_ack_1, ack => convTranspose_CP_39_elements(274)); -- 
    -- CP-element group 275:  transition  input  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	268 
    -- CP-element group 275: successors 
    -- CP-element group 275:  members (3) 
      -- CP-element group 275: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1040_Sample/ra
      -- CP-element group 275: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1040_Sample/$exit
      -- CP-element group 275: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1040_sample_completed_
      -- 
    ra_2186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1040_inst_ack_0, ack => convTranspose_CP_39_elements(275)); -- 
    -- CP-element group 276:  transition  input  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	264 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	296 
    -- CP-element group 276:  members (3) 
      -- CP-element group 276: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1040_Update/ca
      -- CP-element group 276: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1040_Update/$exit
      -- CP-element group 276: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1040_update_completed_
      -- 
    ca_2191_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1040_inst_ack_1, ack => convTranspose_CP_39_elements(276)); -- 
    -- CP-element group 277:  transition  input  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	268 
    -- CP-element group 277: successors 
    -- CP-element group 277:  members (3) 
      -- CP-element group 277: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1050_Sample/ra
      -- CP-element group 277: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1050_Sample/$exit
      -- CP-element group 277: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1050_sample_completed_
      -- 
    ra_2200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1050_inst_ack_0, ack => convTranspose_CP_39_elements(277)); -- 
    -- CP-element group 278:  transition  input  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	264 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	293 
    -- CP-element group 278:  members (3) 
      -- CP-element group 278: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1050_Update/ca
      -- CP-element group 278: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1050_Update/$exit
      -- CP-element group 278: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1050_update_completed_
      -- 
    ca_2205_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1050_inst_ack_1, ack => convTranspose_CP_39_elements(278)); -- 
    -- CP-element group 279:  transition  input  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	268 
    -- CP-element group 279: successors 
    -- CP-element group 279:  members (3) 
      -- CP-element group 279: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1060_Sample/ra
      -- CP-element group 279: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1060_Sample/$exit
      -- CP-element group 279: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1060_sample_completed_
      -- 
    ra_2214_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1060_inst_ack_0, ack => convTranspose_CP_39_elements(279)); -- 
    -- CP-element group 280:  transition  input  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	264 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	290 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1060_Update/$exit
      -- CP-element group 280: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1060_Update/ca
      -- CP-element group 280: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1060_update_completed_
      -- 
    ca_2219_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1060_inst_ack_1, ack => convTranspose_CP_39_elements(280)); -- 
    -- CP-element group 281:  transition  input  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	268 
    -- CP-element group 281: successors 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1070_sample_completed_
      -- CP-element group 281: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1070_Sample/$exit
      -- CP-element group 281: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1070_Sample/ra
      -- 
    ra_2228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1070_inst_ack_0, ack => convTranspose_CP_39_elements(281)); -- 
    -- CP-element group 282:  transition  input  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	264 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	287 
    -- CP-element group 282:  members (3) 
      -- CP-element group 282: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1070_update_completed_
      -- CP-element group 282: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1070_Update/ca
      -- CP-element group 282: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1070_Update/$exit
      -- 
    ca_2233_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1070_inst_ack_1, ack => convTranspose_CP_39_elements(282)); -- 
    -- CP-element group 283:  transition  input  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	268 
    -- CP-element group 283: successors 
    -- CP-element group 283:  members (3) 
      -- CP-element group 283: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1080_Sample/ra
      -- CP-element group 283: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1080_Sample/$exit
      -- CP-element group 283: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1080_sample_completed_
      -- 
    ra_2242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 283_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1080_inst_ack_0, ack => convTranspose_CP_39_elements(283)); -- 
    -- CP-element group 284:  transition  input  output  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	264 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	285 
    -- CP-element group 284:  members (6) 
      -- CP-element group 284: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1082_Sample/$entry
      -- CP-element group 284: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1082_sample_start_
      -- CP-element group 284: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1080_Update/ca
      -- CP-element group 284: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1080_Update/$exit
      -- CP-element group 284: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/type_cast_1080_update_completed_
      -- CP-element group 284: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1082_Sample/req
      -- 
    ca_2247_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1080_inst_ack_1, ack => convTranspose_CP_39_elements(284)); -- 
    req_2255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(284), ack => WPIPE_ConvTranspose_output_pipe_1082_inst_req_0); -- 
    -- CP-element group 285:  transition  input  output  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	284 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	286 
    -- CP-element group 285:  members (6) 
      -- CP-element group 285: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1082_sample_completed_
      -- CP-element group 285: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1082_update_start_
      -- CP-element group 285: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1082_Update/req
      -- CP-element group 285: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1082_Update/$entry
      -- CP-element group 285: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1082_Sample/ack
      -- CP-element group 285: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1082_Sample/$exit
      -- 
    ack_2256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1082_inst_ack_0, ack => convTranspose_CP_39_elements(285)); -- 
    req_2260_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2260_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(285), ack => WPIPE_ConvTranspose_output_pipe_1082_inst_req_1); -- 
    -- CP-element group 286:  transition  input  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	285 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	287 
    -- CP-element group 286:  members (3) 
      -- CP-element group 286: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1082_update_completed_
      -- CP-element group 286: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1082_Update/ack
      -- CP-element group 286: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1082_Update/$exit
      -- 
    ack_2261_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1082_inst_ack_1, ack => convTranspose_CP_39_elements(286)); -- 
    -- CP-element group 287:  join  transition  output  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	282 
    -- CP-element group 287: 	286 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	288 
    -- CP-element group 287:  members (3) 
      -- CP-element group 287: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1085_sample_start_
      -- CP-element group 287: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1085_Sample/$entry
      -- CP-element group 287: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1085_Sample/req
      -- 
    req_2269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(287), ack => WPIPE_ConvTranspose_output_pipe_1085_inst_req_0); -- 
    convTranspose_cp_element_group_287: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_287"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(282) & convTranspose_CP_39_elements(286);
      gj_convTranspose_cp_element_group_287 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(287), clk => clk, reset => reset); --
    end block;
    -- CP-element group 288:  transition  input  output  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	287 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	289 
    -- CP-element group 288:  members (6) 
      -- CP-element group 288: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1085_sample_completed_
      -- CP-element group 288: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1085_update_start_
      -- CP-element group 288: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1085_Sample/$exit
      -- CP-element group 288: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1085_Sample/ack
      -- CP-element group 288: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1085_Update/$entry
      -- CP-element group 288: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1085_Update/req
      -- 
    ack_2270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1085_inst_ack_0, ack => convTranspose_CP_39_elements(288)); -- 
    req_2274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(288), ack => WPIPE_ConvTranspose_output_pipe_1085_inst_req_1); -- 
    -- CP-element group 289:  transition  input  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	288 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	290 
    -- CP-element group 289:  members (3) 
      -- CP-element group 289: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1085_Update/$exit
      -- CP-element group 289: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1085_update_completed_
      -- CP-element group 289: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1085_Update/ack
      -- 
    ack_2275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1085_inst_ack_1, ack => convTranspose_CP_39_elements(289)); -- 
    -- CP-element group 290:  join  transition  output  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	280 
    -- CP-element group 290: 	289 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	291 
    -- CP-element group 290:  members (3) 
      -- CP-element group 290: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1088_Sample/req
      -- CP-element group 290: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1088_sample_start_
      -- CP-element group 290: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1088_Sample/$entry
      -- 
    req_2283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(290), ack => WPIPE_ConvTranspose_output_pipe_1088_inst_req_0); -- 
    convTranspose_cp_element_group_290: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_290"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(280) & convTranspose_CP_39_elements(289);
      gj_convTranspose_cp_element_group_290 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(290), clk => clk, reset => reset); --
    end block;
    -- CP-element group 291:  transition  input  output  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	290 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	292 
    -- CP-element group 291:  members (6) 
      -- CP-element group 291: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1088_Update/req
      -- CP-element group 291: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1088_Update/$entry
      -- CP-element group 291: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1088_Sample/ack
      -- CP-element group 291: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1088_Sample/$exit
      -- CP-element group 291: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1088_update_start_
      -- CP-element group 291: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1088_sample_completed_
      -- 
    ack_2284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1088_inst_ack_0, ack => convTranspose_CP_39_elements(291)); -- 
    req_2288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(291), ack => WPIPE_ConvTranspose_output_pipe_1088_inst_req_1); -- 
    -- CP-element group 292:  transition  input  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	291 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	293 
    -- CP-element group 292:  members (3) 
      -- CP-element group 292: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1088_Update/ack
      -- CP-element group 292: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1088_Update/$exit
      -- CP-element group 292: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1088_update_completed_
      -- 
    ack_2289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1088_inst_ack_1, ack => convTranspose_CP_39_elements(292)); -- 
    -- CP-element group 293:  join  transition  output  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	278 
    -- CP-element group 293: 	292 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	294 
    -- CP-element group 293:  members (3) 
      -- CP-element group 293: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1091_Sample/$entry
      -- CP-element group 293: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1091_Sample/req
      -- CP-element group 293: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1091_sample_start_
      -- 
    req_2297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(293), ack => WPIPE_ConvTranspose_output_pipe_1091_inst_req_0); -- 
    convTranspose_cp_element_group_293: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_293"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(278) & convTranspose_CP_39_elements(292);
      gj_convTranspose_cp_element_group_293 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(293), clk => clk, reset => reset); --
    end block;
    -- CP-element group 294:  transition  input  output  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	293 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	295 
    -- CP-element group 294:  members (6) 
      -- CP-element group 294: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1091_Update/req
      -- CP-element group 294: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1091_Sample/$exit
      -- CP-element group 294: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1091_Sample/ack
      -- CP-element group 294: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1091_Update/$entry
      -- CP-element group 294: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1091_update_start_
      -- CP-element group 294: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1091_sample_completed_
      -- 
    ack_2298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 294_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1091_inst_ack_0, ack => convTranspose_CP_39_elements(294)); -- 
    req_2302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(294), ack => WPIPE_ConvTranspose_output_pipe_1091_inst_req_1); -- 
    -- CP-element group 295:  transition  input  bypass 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	294 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	296 
    -- CP-element group 295:  members (3) 
      -- CP-element group 295: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1091_Update/ack
      -- CP-element group 295: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1091_Update/$exit
      -- CP-element group 295: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1091_update_completed_
      -- 
    ack_2303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1091_inst_ack_1, ack => convTranspose_CP_39_elements(295)); -- 
    -- CP-element group 296:  join  transition  output  bypass 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	276 
    -- CP-element group 296: 	295 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	297 
    -- CP-element group 296:  members (3) 
      -- CP-element group 296: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1094_Sample/$entry
      -- CP-element group 296: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1094_Sample/req
      -- CP-element group 296: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1094_sample_start_
      -- 
    req_2311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(296), ack => WPIPE_ConvTranspose_output_pipe_1094_inst_req_0); -- 
    convTranspose_cp_element_group_296: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_296"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(276) & convTranspose_CP_39_elements(295);
      gj_convTranspose_cp_element_group_296 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(296), clk => clk, reset => reset); --
    end block;
    -- CP-element group 297:  transition  input  output  bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	296 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	298 
    -- CP-element group 297:  members (6) 
      -- CP-element group 297: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1094_Sample/$exit
      -- CP-element group 297: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1094_Sample/ack
      -- CP-element group 297: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1094_Update/$entry
      -- CP-element group 297: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1094_Update/req
      -- CP-element group 297: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1094_update_start_
      -- CP-element group 297: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1094_sample_completed_
      -- 
    ack_2312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1094_inst_ack_0, ack => convTranspose_CP_39_elements(297)); -- 
    req_2316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(297), ack => WPIPE_ConvTranspose_output_pipe_1094_inst_req_1); -- 
    -- CP-element group 298:  transition  input  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	297 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	299 
    -- CP-element group 298:  members (3) 
      -- CP-element group 298: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1094_Update/$exit
      -- CP-element group 298: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1094_update_completed_
      -- CP-element group 298: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1094_Update/ack
      -- 
    ack_2317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 298_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1094_inst_ack_1, ack => convTranspose_CP_39_elements(298)); -- 
    -- CP-element group 299:  join  transition  output  bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	274 
    -- CP-element group 299: 	298 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	300 
    -- CP-element group 299:  members (3) 
      -- CP-element group 299: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1097_Sample/req
      -- CP-element group 299: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1097_Sample/$entry
      -- CP-element group 299: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1097_sample_start_
      -- 
    req_2325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(299), ack => WPIPE_ConvTranspose_output_pipe_1097_inst_req_0); -- 
    convTranspose_cp_element_group_299: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_299"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(274) & convTranspose_CP_39_elements(298);
      gj_convTranspose_cp_element_group_299 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(299), clk => clk, reset => reset); --
    end block;
    -- CP-element group 300:  transition  input  output  bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	299 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	301 
    -- CP-element group 300:  members (6) 
      -- CP-element group 300: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1097_Sample/ack
      -- CP-element group 300: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1097_Update/$entry
      -- CP-element group 300: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1097_Sample/$exit
      -- CP-element group 300: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1097_update_start_
      -- CP-element group 300: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1097_sample_completed_
      -- CP-element group 300: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1097_Update/req
      -- 
    ack_2326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1097_inst_ack_0, ack => convTranspose_CP_39_elements(300)); -- 
    req_2330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(300), ack => WPIPE_ConvTranspose_output_pipe_1097_inst_req_1); -- 
    -- CP-element group 301:  transition  input  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	300 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	302 
    -- CP-element group 301:  members (3) 
      -- CP-element group 301: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1097_Update/$exit
      -- CP-element group 301: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1097_update_completed_
      -- CP-element group 301: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1097_Update/ack
      -- 
    ack_2331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 301_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1097_inst_ack_1, ack => convTranspose_CP_39_elements(301)); -- 
    -- CP-element group 302:  join  transition  output  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	272 
    -- CP-element group 302: 	301 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	303 
    -- CP-element group 302:  members (3) 
      -- CP-element group 302: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1100_Sample/$entry
      -- CP-element group 302: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1100_Sample/req
      -- CP-element group 302: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1100_sample_start_
      -- 
    req_2339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(302), ack => WPIPE_ConvTranspose_output_pipe_1100_inst_req_0); -- 
    convTranspose_cp_element_group_302: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_302"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(272) & convTranspose_CP_39_elements(301);
      gj_convTranspose_cp_element_group_302 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(302), clk => clk, reset => reset); --
    end block;
    -- CP-element group 303:  transition  input  output  bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	302 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	304 
    -- CP-element group 303:  members (6) 
      -- CP-element group 303: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1100_Sample/$exit
      -- CP-element group 303: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1100_update_start_
      -- CP-element group 303: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1100_sample_completed_
      -- CP-element group 303: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1100_Update/req
      -- CP-element group 303: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1100_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1100_Sample/ack
      -- 
    ack_2340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1100_inst_ack_0, ack => convTranspose_CP_39_elements(303)); -- 
    req_2344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(303), ack => WPIPE_ConvTranspose_output_pipe_1100_inst_req_1); -- 
    -- CP-element group 304:  transition  input  bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	303 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	305 
    -- CP-element group 304:  members (3) 
      -- CP-element group 304: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1100_update_completed_
      -- CP-element group 304: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1100_Update/ack
      -- CP-element group 304: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1100_Update/$exit
      -- 
    ack_2345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1100_inst_ack_1, ack => convTranspose_CP_39_elements(304)); -- 
    -- CP-element group 305:  join  transition  output  bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	270 
    -- CP-element group 305: 	304 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	306 
    -- CP-element group 305:  members (3) 
      -- CP-element group 305: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1103_sample_start_
      -- CP-element group 305: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1103_Sample/$entry
      -- CP-element group 305: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1103_Sample/req
      -- 
    req_2353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(305), ack => WPIPE_ConvTranspose_output_pipe_1103_inst_req_0); -- 
    convTranspose_cp_element_group_305: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_305"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(270) & convTranspose_CP_39_elements(304);
      gj_convTranspose_cp_element_group_305 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(305), clk => clk, reset => reset); --
    end block;
    -- CP-element group 306:  transition  input  output  bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	305 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	307 
    -- CP-element group 306:  members (6) 
      -- CP-element group 306: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1103_Update/req
      -- CP-element group 306: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1103_sample_completed_
      -- CP-element group 306: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1103_update_start_
      -- CP-element group 306: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1103_Update/$entry
      -- CP-element group 306: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1103_Sample/ack
      -- CP-element group 306: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1103_Sample/$exit
      -- 
    ack_2354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1103_inst_ack_0, ack => convTranspose_CP_39_elements(306)); -- 
    req_2358_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2358_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(306), ack => WPIPE_ConvTranspose_output_pipe_1103_inst_req_1); -- 
    -- CP-element group 307:  branch  transition  place  input  output  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	306 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	308 
    -- CP-element group 307: 	309 
    -- CP-element group 307:  members (13) 
      -- CP-element group 307: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105__exit__
      -- CP-element group 307: 	 branch_block_stmt_26/if_stmt_1107__entry__
      -- CP-element group 307: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1103_Update/ack
      -- CP-element group 307: 	 branch_block_stmt_26/if_stmt_1107_eval_test/$exit
      -- CP-element group 307: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/$exit
      -- CP-element group 307: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1103_update_completed_
      -- CP-element group 307: 	 branch_block_stmt_26/call_stmt_997_to_assign_stmt_1105/WPIPE_ConvTranspose_output_pipe_1103_Update/$exit
      -- CP-element group 307: 	 branch_block_stmt_26/if_stmt_1107_eval_test/$entry
      -- CP-element group 307: 	 branch_block_stmt_26/if_stmt_1107_else_link/$entry
      -- CP-element group 307: 	 branch_block_stmt_26/if_stmt_1107_dead_link/$entry
      -- CP-element group 307: 	 branch_block_stmt_26/if_stmt_1107_if_link/$entry
      -- CP-element group 307: 	 branch_block_stmt_26/R_cmp264448_1108_place
      -- CP-element group 307: 	 branch_block_stmt_26/if_stmt_1107_eval_test/branch_req
      -- 
    ack_2359_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1103_inst_ack_1, ack => convTranspose_CP_39_elements(307)); -- 
    branch_req_2367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(307), ack => if_stmt_1107_branch_req_0); -- 
    -- CP-element group 308:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	307 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	310 
    -- CP-element group 308: 	311 
    -- CP-element group 308:  members (18) 
      -- CP-element group 308: 	 branch_block_stmt_26/merge_stmt_1113__exit__
      -- CP-element group 308: 	 branch_block_stmt_26/assign_stmt_1119_to_assign_stmt_1148__entry__
      -- CP-element group 308: 	 branch_block_stmt_26/forx_xend273_bbx_xnph
      -- CP-element group 308: 	 branch_block_stmt_26/if_stmt_1107_if_link/if_choice_transition
      -- CP-element group 308: 	 branch_block_stmt_26/if_stmt_1107_if_link/$exit
      -- CP-element group 308: 	 branch_block_stmt_26/assign_stmt_1119_to_assign_stmt_1148/$entry
      -- CP-element group 308: 	 branch_block_stmt_26/assign_stmt_1119_to_assign_stmt_1148/type_cast_1134_sample_start_
      -- CP-element group 308: 	 branch_block_stmt_26/assign_stmt_1119_to_assign_stmt_1148/type_cast_1134_update_start_
      -- CP-element group 308: 	 branch_block_stmt_26/assign_stmt_1119_to_assign_stmt_1148/type_cast_1134_Sample/$entry
      -- CP-element group 308: 	 branch_block_stmt_26/assign_stmt_1119_to_assign_stmt_1148/type_cast_1134_Sample/rr
      -- CP-element group 308: 	 branch_block_stmt_26/assign_stmt_1119_to_assign_stmt_1148/type_cast_1134_Update/$entry
      -- CP-element group 308: 	 branch_block_stmt_26/assign_stmt_1119_to_assign_stmt_1148/type_cast_1134_Update/cr
      -- CP-element group 308: 	 branch_block_stmt_26/forx_xend273_bbx_xnph_PhiReq/$entry
      -- CP-element group 308: 	 branch_block_stmt_26/forx_xend273_bbx_xnph_PhiReq/$exit
      -- CP-element group 308: 	 branch_block_stmt_26/merge_stmt_1113_PhiReqMerge
      -- CP-element group 308: 	 branch_block_stmt_26/merge_stmt_1113_PhiAck/$entry
      -- CP-element group 308: 	 branch_block_stmt_26/merge_stmt_1113_PhiAck/$exit
      -- CP-element group 308: 	 branch_block_stmt_26/merge_stmt_1113_PhiAck/dummy
      -- 
    if_choice_transition_2372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1107_branch_ack_1, ack => convTranspose_CP_39_elements(308)); -- 
    rr_2389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(308), ack => type_cast_1134_inst_req_0); -- 
    cr_2394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(308), ack => type_cast_1134_inst_req_1); -- 
    -- CP-element group 309:  transition  place  input  bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	307 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	387 
    -- CP-element group 309:  members (5) 
      -- CP-element group 309: 	 branch_block_stmt_26/forx_xend273_forx_xend443_PhiReq/$exit
      -- CP-element group 309: 	 branch_block_stmt_26/if_stmt_1107_else_link/else_choice_transition
      -- CP-element group 309: 	 branch_block_stmt_26/if_stmt_1107_else_link/$exit
      -- CP-element group 309: 	 branch_block_stmt_26/forx_xend273_forx_xend443_PhiReq/$entry
      -- CP-element group 309: 	 branch_block_stmt_26/forx_xend273_forx_xend443
      -- 
    else_choice_transition_2376_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 309_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1107_branch_ack_0, ack => convTranspose_CP_39_elements(309)); -- 
    -- CP-element group 310:  transition  input  bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	308 
    -- CP-element group 310: successors 
    -- CP-element group 310:  members (3) 
      -- CP-element group 310: 	 branch_block_stmt_26/assign_stmt_1119_to_assign_stmt_1148/type_cast_1134_sample_completed_
      -- CP-element group 310: 	 branch_block_stmt_26/assign_stmt_1119_to_assign_stmt_1148/type_cast_1134_Sample/$exit
      -- CP-element group 310: 	 branch_block_stmt_26/assign_stmt_1119_to_assign_stmt_1148/type_cast_1134_Sample/ra
      -- 
    ra_2390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 310_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1134_inst_ack_0, ack => convTranspose_CP_39_elements(310)); -- 
    -- CP-element group 311:  transition  place  input  bypass 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	308 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	381 
    -- CP-element group 311:  members (9) 
      -- CP-element group 311: 	 branch_block_stmt_26/assign_stmt_1119_to_assign_stmt_1148__exit__
      -- CP-element group 311: 	 branch_block_stmt_26/bbx_xnph_forx_xbody370
      -- CP-element group 311: 	 branch_block_stmt_26/assign_stmt_1119_to_assign_stmt_1148/$exit
      -- CP-element group 311: 	 branch_block_stmt_26/assign_stmt_1119_to_assign_stmt_1148/type_cast_1134_update_completed_
      -- CP-element group 311: 	 branch_block_stmt_26/assign_stmt_1119_to_assign_stmt_1148/type_cast_1134_Update/$exit
      -- CP-element group 311: 	 branch_block_stmt_26/assign_stmt_1119_to_assign_stmt_1148/type_cast_1134_Update/ca
      -- CP-element group 311: 	 branch_block_stmt_26/bbx_xnph_forx_xbody370_PhiReq/$entry
      -- CP-element group 311: 	 branch_block_stmt_26/bbx_xnph_forx_xbody370_PhiReq/phi_stmt_1151/$entry
      -- CP-element group 311: 	 branch_block_stmt_26/bbx_xnph_forx_xbody370_PhiReq/phi_stmt_1151/phi_stmt_1151_sources/$entry
      -- 
    ca_2395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1134_inst_ack_1, ack => convTranspose_CP_39_elements(311)); -- 
    -- CP-element group 312:  transition  input  bypass 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	386 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	357 
    -- CP-element group 312:  members (3) 
      -- CP-element group 312: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/array_obj_ref_1163_final_index_sum_regn_sample_complete
      -- CP-element group 312: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/array_obj_ref_1163_final_index_sum_regn_Sample/$exit
      -- CP-element group 312: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/array_obj_ref_1163_final_index_sum_regn_Sample/ack
      -- 
    ack_2424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1163_index_offset_ack_0, ack => convTranspose_CP_39_elements(312)); -- 
    -- CP-element group 313:  transition  input  output  bypass 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	386 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	314 
    -- CP-element group 313:  members (11) 
      -- CP-element group 313: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/addr_of_1164_sample_start_
      -- CP-element group 313: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/array_obj_ref_1163_root_address_calculated
      -- CP-element group 313: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/array_obj_ref_1163_offset_calculated
      -- CP-element group 313: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/array_obj_ref_1163_final_index_sum_regn_Update/$exit
      -- CP-element group 313: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/array_obj_ref_1163_final_index_sum_regn_Update/ack
      -- CP-element group 313: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/array_obj_ref_1163_base_plus_offset/$entry
      -- CP-element group 313: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/array_obj_ref_1163_base_plus_offset/$exit
      -- CP-element group 313: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/array_obj_ref_1163_base_plus_offset/sum_rename_req
      -- CP-element group 313: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/array_obj_ref_1163_base_plus_offset/sum_rename_ack
      -- CP-element group 313: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/addr_of_1164_request/$entry
      -- CP-element group 313: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/addr_of_1164_request/req
      -- 
    ack_2429_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1163_index_offset_ack_1, ack => convTranspose_CP_39_elements(313)); -- 
    req_2438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(313), ack => addr_of_1164_final_reg_req_0); -- 
    -- CP-element group 314:  transition  input  bypass 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	313 
    -- CP-element group 314: successors 
    -- CP-element group 314:  members (3) 
      -- CP-element group 314: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/addr_of_1164_sample_completed_
      -- CP-element group 314: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/addr_of_1164_request/$exit
      -- CP-element group 314: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/addr_of_1164_request/ack
      -- 
    ack_2439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1164_final_reg_ack_0, ack => convTranspose_CP_39_elements(314)); -- 
    -- CP-element group 315:  join  fork  transition  input  output  bypass 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	386 
    -- CP-element group 315: successors 
    -- CP-element group 315: 	316 
    -- CP-element group 315:  members (24) 
      -- CP-element group 315: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/addr_of_1164_update_completed_
      -- CP-element group 315: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/addr_of_1164_complete/$exit
      -- CP-element group 315: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/addr_of_1164_complete/ack
      -- CP-element group 315: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/ptr_deref_1168_sample_start_
      -- CP-element group 315: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/ptr_deref_1168_base_address_calculated
      -- CP-element group 315: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/ptr_deref_1168_word_address_calculated
      -- CP-element group 315: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/ptr_deref_1168_root_address_calculated
      -- CP-element group 315: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/ptr_deref_1168_base_address_resized
      -- CP-element group 315: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/ptr_deref_1168_base_addr_resize/$entry
      -- CP-element group 315: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/ptr_deref_1168_base_addr_resize/$exit
      -- CP-element group 315: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/ptr_deref_1168_base_addr_resize/base_resize_req
      -- CP-element group 315: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/ptr_deref_1168_base_addr_resize/base_resize_ack
      -- CP-element group 315: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/ptr_deref_1168_base_plus_offset/$entry
      -- CP-element group 315: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/ptr_deref_1168_base_plus_offset/$exit
      -- CP-element group 315: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/ptr_deref_1168_base_plus_offset/sum_rename_req
      -- CP-element group 315: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/ptr_deref_1168_base_plus_offset/sum_rename_ack
      -- CP-element group 315: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/ptr_deref_1168_word_addrgen/$entry
      -- CP-element group 315: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/ptr_deref_1168_word_addrgen/$exit
      -- CP-element group 315: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/ptr_deref_1168_word_addrgen/root_register_req
      -- CP-element group 315: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/ptr_deref_1168_word_addrgen/root_register_ack
      -- CP-element group 315: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/ptr_deref_1168_Sample/$entry
      -- CP-element group 315: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/ptr_deref_1168_Sample/word_access_start/$entry
      -- CP-element group 315: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/ptr_deref_1168_Sample/word_access_start/word_0/$entry
      -- CP-element group 315: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/ptr_deref_1168_Sample/word_access_start/word_0/rr
      -- 
    ack_2444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1164_final_reg_ack_1, ack => convTranspose_CP_39_elements(315)); -- 
    rr_2477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(315), ack => ptr_deref_1168_load_0_req_0); -- 
    -- CP-element group 316:  transition  input  bypass 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	315 
    -- CP-element group 316: successors 
    -- CP-element group 316:  members (5) 
      -- CP-element group 316: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/ptr_deref_1168_sample_completed_
      -- CP-element group 316: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/ptr_deref_1168_Sample/$exit
      -- CP-element group 316: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/ptr_deref_1168_Sample/word_access_start/$exit
      -- CP-element group 316: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/ptr_deref_1168_Sample/word_access_start/word_0/$exit
      -- CP-element group 316: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/ptr_deref_1168_Sample/word_access_start/word_0/ra
      -- 
    ra_2478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1168_load_0_ack_0, ack => convTranspose_CP_39_elements(316)); -- 
    -- CP-element group 317:  fork  transition  input  output  bypass 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	386 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	318 
    -- CP-element group 317: 	320 
    -- CP-element group 317: 	322 
    -- CP-element group 317: 	324 
    -- CP-element group 317: 	326 
    -- CP-element group 317: 	328 
    -- CP-element group 317: 	330 
    -- CP-element group 317: 	332 
    -- CP-element group 317:  members (33) 
      -- CP-element group 317: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/ptr_deref_1168_update_completed_
      -- CP-element group 317: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/ptr_deref_1168_Update/$exit
      -- CP-element group 317: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/ptr_deref_1168_Update/word_access_complete/$exit
      -- CP-element group 317: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/ptr_deref_1168_Update/word_access_complete/word_0/$exit
      -- CP-element group 317: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/ptr_deref_1168_Update/word_access_complete/word_0/ca
      -- CP-element group 317: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/ptr_deref_1168_Update/ptr_deref_1168_Merge/$entry
      -- CP-element group 317: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/ptr_deref_1168_Update/ptr_deref_1168_Merge/$exit
      -- CP-element group 317: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/ptr_deref_1168_Update/ptr_deref_1168_Merge/merge_req
      -- CP-element group 317: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/ptr_deref_1168_Update/ptr_deref_1168_Merge/merge_ack
      -- CP-element group 317: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1172_sample_start_
      -- CP-element group 317: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1172_Sample/$entry
      -- CP-element group 317: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1172_Sample/rr
      -- CP-element group 317: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1182_sample_start_
      -- CP-element group 317: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1182_Sample/$entry
      -- CP-element group 317: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1182_Sample/rr
      -- CP-element group 317: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1192_sample_start_
      -- CP-element group 317: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1192_Sample/$entry
      -- CP-element group 317: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1192_Sample/rr
      -- CP-element group 317: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1202_sample_start_
      -- CP-element group 317: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1202_Sample/$entry
      -- CP-element group 317: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1202_Sample/rr
      -- CP-element group 317: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1212_sample_start_
      -- CP-element group 317: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1212_Sample/$entry
      -- CP-element group 317: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1212_Sample/rr
      -- CP-element group 317: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1222_sample_start_
      -- CP-element group 317: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1222_Sample/$entry
      -- CP-element group 317: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1222_Sample/rr
      -- CP-element group 317: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1232_sample_start_
      -- CP-element group 317: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1232_Sample/$entry
      -- CP-element group 317: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1232_Sample/rr
      -- CP-element group 317: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1242_sample_start_
      -- CP-element group 317: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1242_Sample/$entry
      -- CP-element group 317: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1242_Sample/rr
      -- 
    ca_2489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 317_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1168_load_0_ack_1, ack => convTranspose_CP_39_elements(317)); -- 
    rr_2502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(317), ack => type_cast_1172_inst_req_0); -- 
    rr_2516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(317), ack => type_cast_1182_inst_req_0); -- 
    rr_2530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(317), ack => type_cast_1192_inst_req_0); -- 
    rr_2544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(317), ack => type_cast_1202_inst_req_0); -- 
    rr_2558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(317), ack => type_cast_1212_inst_req_0); -- 
    rr_2572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(317), ack => type_cast_1222_inst_req_0); -- 
    rr_2586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(317), ack => type_cast_1232_inst_req_0); -- 
    rr_2600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(317), ack => type_cast_1242_inst_req_0); -- 
    -- CP-element group 318:  transition  input  bypass 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	317 
    -- CP-element group 318: successors 
    -- CP-element group 318:  members (3) 
      -- CP-element group 318: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1172_sample_completed_
      -- CP-element group 318: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1172_Sample/$exit
      -- CP-element group 318: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1172_Sample/ra
      -- 
    ra_2503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 318_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1172_inst_ack_0, ack => convTranspose_CP_39_elements(318)); -- 
    -- CP-element group 319:  transition  input  bypass 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	386 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	354 
    -- CP-element group 319:  members (3) 
      -- CP-element group 319: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1172_update_completed_
      -- CP-element group 319: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1172_Update/$exit
      -- CP-element group 319: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1172_Update/ca
      -- 
    ca_2508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 319_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1172_inst_ack_1, ack => convTranspose_CP_39_elements(319)); -- 
    -- CP-element group 320:  transition  input  bypass 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	317 
    -- CP-element group 320: successors 
    -- CP-element group 320:  members (3) 
      -- CP-element group 320: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1182_sample_completed_
      -- CP-element group 320: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1182_Sample/$exit
      -- CP-element group 320: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1182_Sample/ra
      -- 
    ra_2517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 320_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1182_inst_ack_0, ack => convTranspose_CP_39_elements(320)); -- 
    -- CP-element group 321:  transition  input  bypass 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	386 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	351 
    -- CP-element group 321:  members (3) 
      -- CP-element group 321: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1182_update_completed_
      -- CP-element group 321: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1182_Update/$exit
      -- CP-element group 321: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1182_Update/ca
      -- 
    ca_2522_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1182_inst_ack_1, ack => convTranspose_CP_39_elements(321)); -- 
    -- CP-element group 322:  transition  input  bypass 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	317 
    -- CP-element group 322: successors 
    -- CP-element group 322:  members (3) 
      -- CP-element group 322: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1192_sample_completed_
      -- CP-element group 322: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1192_Sample/$exit
      -- CP-element group 322: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1192_Sample/ra
      -- 
    ra_2531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 322_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1192_inst_ack_0, ack => convTranspose_CP_39_elements(322)); -- 
    -- CP-element group 323:  transition  input  bypass 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	386 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	348 
    -- CP-element group 323:  members (3) 
      -- CP-element group 323: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1192_update_completed_
      -- CP-element group 323: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1192_Update/$exit
      -- CP-element group 323: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1192_Update/ca
      -- 
    ca_2536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 323_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1192_inst_ack_1, ack => convTranspose_CP_39_elements(323)); -- 
    -- CP-element group 324:  transition  input  bypass 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	317 
    -- CP-element group 324: successors 
    -- CP-element group 324:  members (3) 
      -- CP-element group 324: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1202_sample_completed_
      -- CP-element group 324: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1202_Sample/$exit
      -- CP-element group 324: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1202_Sample/ra
      -- 
    ra_2545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 324_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1202_inst_ack_0, ack => convTranspose_CP_39_elements(324)); -- 
    -- CP-element group 325:  transition  input  bypass 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	386 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	345 
    -- CP-element group 325:  members (3) 
      -- CP-element group 325: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1202_update_completed_
      -- CP-element group 325: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1202_Update/$exit
      -- CP-element group 325: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1202_Update/ca
      -- 
    ca_2550_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 325_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1202_inst_ack_1, ack => convTranspose_CP_39_elements(325)); -- 
    -- CP-element group 326:  transition  input  bypass 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	317 
    -- CP-element group 326: successors 
    -- CP-element group 326:  members (3) 
      -- CP-element group 326: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1212_sample_completed_
      -- CP-element group 326: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1212_Sample/$exit
      -- CP-element group 326: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1212_Sample/ra
      -- 
    ra_2559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 326_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1212_inst_ack_0, ack => convTranspose_CP_39_elements(326)); -- 
    -- CP-element group 327:  transition  input  bypass 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	386 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	342 
    -- CP-element group 327:  members (3) 
      -- CP-element group 327: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1212_update_completed_
      -- CP-element group 327: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1212_Update/$exit
      -- CP-element group 327: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1212_Update/ca
      -- 
    ca_2564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 327_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1212_inst_ack_1, ack => convTranspose_CP_39_elements(327)); -- 
    -- CP-element group 328:  transition  input  bypass 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	317 
    -- CP-element group 328: successors 
    -- CP-element group 328:  members (3) 
      -- CP-element group 328: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1222_sample_completed_
      -- CP-element group 328: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1222_Sample/$exit
      -- CP-element group 328: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1222_Sample/ra
      -- 
    ra_2573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 328_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1222_inst_ack_0, ack => convTranspose_CP_39_elements(328)); -- 
    -- CP-element group 329:  transition  input  bypass 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	386 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	339 
    -- CP-element group 329:  members (3) 
      -- CP-element group 329: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1222_update_completed_
      -- CP-element group 329: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1222_Update/$exit
      -- CP-element group 329: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1222_Update/ca
      -- 
    ca_2578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 329_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1222_inst_ack_1, ack => convTranspose_CP_39_elements(329)); -- 
    -- CP-element group 330:  transition  input  bypass 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	317 
    -- CP-element group 330: successors 
    -- CP-element group 330:  members (3) 
      -- CP-element group 330: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1232_sample_completed_
      -- CP-element group 330: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1232_Sample/$exit
      -- CP-element group 330: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1232_Sample/ra
      -- 
    ra_2587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 330_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1232_inst_ack_0, ack => convTranspose_CP_39_elements(330)); -- 
    -- CP-element group 331:  transition  input  bypass 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	386 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	336 
    -- CP-element group 331:  members (3) 
      -- CP-element group 331: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1232_update_completed_
      -- CP-element group 331: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1232_Update/$exit
      -- CP-element group 331: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1232_Update/ca
      -- 
    ca_2592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 331_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1232_inst_ack_1, ack => convTranspose_CP_39_elements(331)); -- 
    -- CP-element group 332:  transition  input  bypass 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	317 
    -- CP-element group 332: successors 
    -- CP-element group 332:  members (3) 
      -- CP-element group 332: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1242_sample_completed_
      -- CP-element group 332: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1242_Sample/$exit
      -- CP-element group 332: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1242_Sample/ra
      -- 
    ra_2601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1242_inst_ack_0, ack => convTranspose_CP_39_elements(332)); -- 
    -- CP-element group 333:  transition  input  output  bypass 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	386 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	334 
    -- CP-element group 333:  members (6) 
      -- CP-element group 333: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1242_update_completed_
      -- CP-element group 333: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1242_Update/$exit
      -- CP-element group 333: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1242_Update/ca
      -- CP-element group 333: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1244_sample_start_
      -- CP-element group 333: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1244_Sample/$entry
      -- CP-element group 333: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1244_Sample/req
      -- 
    ca_2606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 333_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1242_inst_ack_1, ack => convTranspose_CP_39_elements(333)); -- 
    req_2614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(333), ack => WPIPE_ConvTranspose_output_pipe_1244_inst_req_0); -- 
    -- CP-element group 334:  transition  input  output  bypass 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	333 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	335 
    -- CP-element group 334:  members (6) 
      -- CP-element group 334: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1244_sample_completed_
      -- CP-element group 334: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1244_update_start_
      -- CP-element group 334: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1244_Sample/$exit
      -- CP-element group 334: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1244_Sample/ack
      -- CP-element group 334: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1244_Update/$entry
      -- CP-element group 334: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1244_Update/req
      -- 
    ack_2615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 334_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1244_inst_ack_0, ack => convTranspose_CP_39_elements(334)); -- 
    req_2619_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2619_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(334), ack => WPIPE_ConvTranspose_output_pipe_1244_inst_req_1); -- 
    -- CP-element group 335:  transition  input  bypass 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	334 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	336 
    -- CP-element group 335:  members (3) 
      -- CP-element group 335: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1244_update_completed_
      -- CP-element group 335: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1244_Update/$exit
      -- CP-element group 335: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1244_Update/ack
      -- 
    ack_2620_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 335_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1244_inst_ack_1, ack => convTranspose_CP_39_elements(335)); -- 
    -- CP-element group 336:  join  transition  output  bypass 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	331 
    -- CP-element group 336: 	335 
    -- CP-element group 336: successors 
    -- CP-element group 336: 	337 
    -- CP-element group 336:  members (3) 
      -- CP-element group 336: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1247_sample_start_
      -- CP-element group 336: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1247_Sample/$entry
      -- CP-element group 336: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1247_Sample/req
      -- 
    req_2628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(336), ack => WPIPE_ConvTranspose_output_pipe_1247_inst_req_0); -- 
    convTranspose_cp_element_group_336: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_336"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(331) & convTranspose_CP_39_elements(335);
      gj_convTranspose_cp_element_group_336 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(336), clk => clk, reset => reset); --
    end block;
    -- CP-element group 337:  transition  input  output  bypass 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	336 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	338 
    -- CP-element group 337:  members (6) 
      -- CP-element group 337: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1247_sample_completed_
      -- CP-element group 337: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1247_update_start_
      -- CP-element group 337: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1247_Sample/$exit
      -- CP-element group 337: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1247_Sample/ack
      -- CP-element group 337: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1247_Update/$entry
      -- CP-element group 337: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1247_Update/req
      -- 
    ack_2629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1247_inst_ack_0, ack => convTranspose_CP_39_elements(337)); -- 
    req_2633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(337), ack => WPIPE_ConvTranspose_output_pipe_1247_inst_req_1); -- 
    -- CP-element group 338:  transition  input  bypass 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	337 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	339 
    -- CP-element group 338:  members (3) 
      -- CP-element group 338: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1247_update_completed_
      -- CP-element group 338: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1247_Update/$exit
      -- CP-element group 338: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1247_Update/ack
      -- 
    ack_2634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 338_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1247_inst_ack_1, ack => convTranspose_CP_39_elements(338)); -- 
    -- CP-element group 339:  join  transition  output  bypass 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	329 
    -- CP-element group 339: 	338 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	340 
    -- CP-element group 339:  members (3) 
      -- CP-element group 339: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1250_sample_start_
      -- CP-element group 339: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1250_Sample/$entry
      -- CP-element group 339: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1250_Sample/req
      -- 
    req_2642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(339), ack => WPIPE_ConvTranspose_output_pipe_1250_inst_req_0); -- 
    convTranspose_cp_element_group_339: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_339"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(329) & convTranspose_CP_39_elements(338);
      gj_convTranspose_cp_element_group_339 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(339), clk => clk, reset => reset); --
    end block;
    -- CP-element group 340:  transition  input  output  bypass 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	339 
    -- CP-element group 340: successors 
    -- CP-element group 340: 	341 
    -- CP-element group 340:  members (6) 
      -- CP-element group 340: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1250_sample_completed_
      -- CP-element group 340: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1250_update_start_
      -- CP-element group 340: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1250_Sample/$exit
      -- CP-element group 340: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1250_Sample/ack
      -- CP-element group 340: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1250_Update/$entry
      -- CP-element group 340: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1250_Update/req
      -- 
    ack_2643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1250_inst_ack_0, ack => convTranspose_CP_39_elements(340)); -- 
    req_2647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(340), ack => WPIPE_ConvTranspose_output_pipe_1250_inst_req_1); -- 
    -- CP-element group 341:  transition  input  bypass 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	340 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	342 
    -- CP-element group 341:  members (3) 
      -- CP-element group 341: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1250_update_completed_
      -- CP-element group 341: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1250_Update/$exit
      -- CP-element group 341: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1250_Update/ack
      -- 
    ack_2648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1250_inst_ack_1, ack => convTranspose_CP_39_elements(341)); -- 
    -- CP-element group 342:  join  transition  output  bypass 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	327 
    -- CP-element group 342: 	341 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	343 
    -- CP-element group 342:  members (3) 
      -- CP-element group 342: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1253_sample_start_
      -- CP-element group 342: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1253_Sample/$entry
      -- CP-element group 342: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1253_Sample/req
      -- 
    req_2656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(342), ack => WPIPE_ConvTranspose_output_pipe_1253_inst_req_0); -- 
    convTranspose_cp_element_group_342: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_342"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(327) & convTranspose_CP_39_elements(341);
      gj_convTranspose_cp_element_group_342 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(342), clk => clk, reset => reset); --
    end block;
    -- CP-element group 343:  transition  input  output  bypass 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	342 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	344 
    -- CP-element group 343:  members (6) 
      -- CP-element group 343: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1253_sample_completed_
      -- CP-element group 343: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1253_update_start_
      -- CP-element group 343: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1253_Sample/$exit
      -- CP-element group 343: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1253_Sample/ack
      -- CP-element group 343: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1253_Update/$entry
      -- CP-element group 343: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1253_Update/req
      -- 
    ack_2657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 343_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1253_inst_ack_0, ack => convTranspose_CP_39_elements(343)); -- 
    req_2661_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2661_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(343), ack => WPIPE_ConvTranspose_output_pipe_1253_inst_req_1); -- 
    -- CP-element group 344:  transition  input  bypass 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	343 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	345 
    -- CP-element group 344:  members (3) 
      -- CP-element group 344: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1253_update_completed_
      -- CP-element group 344: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1253_Update/$exit
      -- CP-element group 344: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1253_Update/ack
      -- 
    ack_2662_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 344_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1253_inst_ack_1, ack => convTranspose_CP_39_elements(344)); -- 
    -- CP-element group 345:  join  transition  output  bypass 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	325 
    -- CP-element group 345: 	344 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	346 
    -- CP-element group 345:  members (3) 
      -- CP-element group 345: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1256_sample_start_
      -- CP-element group 345: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1256_Sample/$entry
      -- CP-element group 345: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1256_Sample/req
      -- 
    req_2670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(345), ack => WPIPE_ConvTranspose_output_pipe_1256_inst_req_0); -- 
    convTranspose_cp_element_group_345: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_345"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(325) & convTranspose_CP_39_elements(344);
      gj_convTranspose_cp_element_group_345 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(345), clk => clk, reset => reset); --
    end block;
    -- CP-element group 346:  transition  input  output  bypass 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	345 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	347 
    -- CP-element group 346:  members (6) 
      -- CP-element group 346: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1256_sample_completed_
      -- CP-element group 346: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1256_update_start_
      -- CP-element group 346: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1256_Sample/$exit
      -- CP-element group 346: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1256_Sample/ack
      -- CP-element group 346: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1256_Update/$entry
      -- CP-element group 346: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1256_Update/req
      -- 
    ack_2671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 346_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1256_inst_ack_0, ack => convTranspose_CP_39_elements(346)); -- 
    req_2675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(346), ack => WPIPE_ConvTranspose_output_pipe_1256_inst_req_1); -- 
    -- CP-element group 347:  transition  input  bypass 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	346 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	348 
    -- CP-element group 347:  members (3) 
      -- CP-element group 347: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1256_update_completed_
      -- CP-element group 347: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1256_Update/$exit
      -- CP-element group 347: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1256_Update/ack
      -- 
    ack_2676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 347_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1256_inst_ack_1, ack => convTranspose_CP_39_elements(347)); -- 
    -- CP-element group 348:  join  transition  output  bypass 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	323 
    -- CP-element group 348: 	347 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	349 
    -- CP-element group 348:  members (3) 
      -- CP-element group 348: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1259_sample_start_
      -- CP-element group 348: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1259_Sample/$entry
      -- CP-element group 348: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1259_Sample/req
      -- 
    req_2684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(348), ack => WPIPE_ConvTranspose_output_pipe_1259_inst_req_0); -- 
    convTranspose_cp_element_group_348: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_348"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(323) & convTranspose_CP_39_elements(347);
      gj_convTranspose_cp_element_group_348 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(348), clk => clk, reset => reset); --
    end block;
    -- CP-element group 349:  transition  input  output  bypass 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	348 
    -- CP-element group 349: successors 
    -- CP-element group 349: 	350 
    -- CP-element group 349:  members (6) 
      -- CP-element group 349: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1259_sample_completed_
      -- CP-element group 349: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1259_update_start_
      -- CP-element group 349: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1259_Sample/$exit
      -- CP-element group 349: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1259_Sample/ack
      -- CP-element group 349: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1259_Update/$entry
      -- CP-element group 349: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1259_Update/req
      -- 
    ack_2685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 349_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1259_inst_ack_0, ack => convTranspose_CP_39_elements(349)); -- 
    req_2689_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2689_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(349), ack => WPIPE_ConvTranspose_output_pipe_1259_inst_req_1); -- 
    -- CP-element group 350:  transition  input  bypass 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	349 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	351 
    -- CP-element group 350:  members (3) 
      -- CP-element group 350: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1259_update_completed_
      -- CP-element group 350: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1259_Update/$exit
      -- CP-element group 350: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1259_Update/ack
      -- 
    ack_2690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 350_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1259_inst_ack_1, ack => convTranspose_CP_39_elements(350)); -- 
    -- CP-element group 351:  join  transition  output  bypass 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	321 
    -- CP-element group 351: 	350 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	352 
    -- CP-element group 351:  members (3) 
      -- CP-element group 351: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1262_sample_start_
      -- CP-element group 351: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1262_Sample/$entry
      -- CP-element group 351: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1262_Sample/req
      -- 
    req_2698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(351), ack => WPIPE_ConvTranspose_output_pipe_1262_inst_req_0); -- 
    convTranspose_cp_element_group_351: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_351"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(321) & convTranspose_CP_39_elements(350);
      gj_convTranspose_cp_element_group_351 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(351), clk => clk, reset => reset); --
    end block;
    -- CP-element group 352:  transition  input  output  bypass 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	351 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	353 
    -- CP-element group 352:  members (6) 
      -- CP-element group 352: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1262_sample_completed_
      -- CP-element group 352: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1262_update_start_
      -- CP-element group 352: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1262_Sample/$exit
      -- CP-element group 352: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1262_Sample/ack
      -- CP-element group 352: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1262_Update/$entry
      -- CP-element group 352: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1262_Update/req
      -- 
    ack_2699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1262_inst_ack_0, ack => convTranspose_CP_39_elements(352)); -- 
    req_2703_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2703_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(352), ack => WPIPE_ConvTranspose_output_pipe_1262_inst_req_1); -- 
    -- CP-element group 353:  transition  input  bypass 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	352 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	354 
    -- CP-element group 353:  members (3) 
      -- CP-element group 353: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1262_update_completed_
      -- CP-element group 353: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1262_Update/$exit
      -- CP-element group 353: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1262_Update/ack
      -- 
    ack_2704_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 353_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1262_inst_ack_1, ack => convTranspose_CP_39_elements(353)); -- 
    -- CP-element group 354:  join  transition  output  bypass 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	319 
    -- CP-element group 354: 	353 
    -- CP-element group 354: successors 
    -- CP-element group 354: 	355 
    -- CP-element group 354:  members (3) 
      -- CP-element group 354: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1265_sample_start_
      -- CP-element group 354: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1265_Sample/$entry
      -- CP-element group 354: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1265_Sample/req
      -- 
    req_2712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(354), ack => WPIPE_ConvTranspose_output_pipe_1265_inst_req_0); -- 
    convTranspose_cp_element_group_354: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_354"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(319) & convTranspose_CP_39_elements(353);
      gj_convTranspose_cp_element_group_354 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(354), clk => clk, reset => reset); --
    end block;
    -- CP-element group 355:  transition  input  output  bypass 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	354 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	356 
    -- CP-element group 355:  members (6) 
      -- CP-element group 355: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1265_sample_completed_
      -- CP-element group 355: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1265_update_start_
      -- CP-element group 355: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1265_Sample/$exit
      -- CP-element group 355: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1265_Sample/ack
      -- CP-element group 355: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1265_Update/$entry
      -- CP-element group 355: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1265_Update/req
      -- 
    ack_2713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 355_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1265_inst_ack_0, ack => convTranspose_CP_39_elements(355)); -- 
    req_2717_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2717_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(355), ack => WPIPE_ConvTranspose_output_pipe_1265_inst_req_1); -- 
    -- CP-element group 356:  transition  input  bypass 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	355 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	357 
    -- CP-element group 356:  members (3) 
      -- CP-element group 356: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1265_update_completed_
      -- CP-element group 356: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1265_Update/$exit
      -- CP-element group 356: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/WPIPE_ConvTranspose_output_pipe_1265_Update/ack
      -- 
    ack_2718_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 356_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1265_inst_ack_1, ack => convTranspose_CP_39_elements(356)); -- 
    -- CP-element group 357:  branch  join  transition  place  output  bypass 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	312 
    -- CP-element group 357: 	356 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	358 
    -- CP-element group 357: 	359 
    -- CP-element group 357:  members (10) 
      -- CP-element group 357: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278__exit__
      -- CP-element group 357: 	 branch_block_stmt_26/if_stmt_1279__entry__
      -- CP-element group 357: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/$exit
      -- CP-element group 357: 	 branch_block_stmt_26/if_stmt_1279_dead_link/$entry
      -- CP-element group 357: 	 branch_block_stmt_26/if_stmt_1279_eval_test/$entry
      -- CP-element group 357: 	 branch_block_stmt_26/if_stmt_1279_eval_test/$exit
      -- CP-element group 357: 	 branch_block_stmt_26/if_stmt_1279_eval_test/branch_req
      -- CP-element group 357: 	 branch_block_stmt_26/R_exitcond1_1280_place
      -- CP-element group 357: 	 branch_block_stmt_26/if_stmt_1279_if_link/$entry
      -- CP-element group 357: 	 branch_block_stmt_26/if_stmt_1279_else_link/$entry
      -- 
    branch_req_2726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(357), ack => if_stmt_1279_branch_req_0); -- 
    convTranspose_cp_element_group_357: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_357"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(312) & convTranspose_CP_39_elements(356);
      gj_convTranspose_cp_element_group_357 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(357), clk => clk, reset => reset); --
    end block;
    -- CP-element group 358:  merge  transition  place  input  bypass 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	357 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	387 
    -- CP-element group 358:  members (13) 
      -- CP-element group 358: 	 branch_block_stmt_26/merge_stmt_1285__exit__
      -- CP-element group 358: 	 branch_block_stmt_26/forx_xend443x_xloopexit_forx_xend443
      -- CP-element group 358: 	 branch_block_stmt_26/forx_xend443x_xloopexit_forx_xend443_PhiReq/$entry
      -- CP-element group 358: 	 branch_block_stmt_26/merge_stmt_1285_PhiAck/dummy
      -- CP-element group 358: 	 branch_block_stmt_26/merge_stmt_1285_PhiAck/$entry
      -- CP-element group 358: 	 branch_block_stmt_26/merge_stmt_1285_PhiAck/$exit
      -- CP-element group 358: 	 branch_block_stmt_26/forx_xbody370_forx_xend443x_xloopexit_PhiReq/$exit
      -- CP-element group 358: 	 branch_block_stmt_26/forx_xbody370_forx_xend443x_xloopexit_PhiReq/$entry
      -- CP-element group 358: 	 branch_block_stmt_26/if_stmt_1279_if_link/$exit
      -- CP-element group 358: 	 branch_block_stmt_26/if_stmt_1279_if_link/if_choice_transition
      -- CP-element group 358: 	 branch_block_stmt_26/forx_xend443x_xloopexit_forx_xend443_PhiReq/$exit
      -- CP-element group 358: 	 branch_block_stmt_26/forx_xbody370_forx_xend443x_xloopexit
      -- CP-element group 358: 	 branch_block_stmt_26/merge_stmt_1285_PhiReqMerge
      -- 
    if_choice_transition_2731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 358_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1279_branch_ack_1, ack => convTranspose_CP_39_elements(358)); -- 
    -- CP-element group 359:  fork  transition  place  input  output  bypass 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	357 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	382 
    -- CP-element group 359: 	383 
    -- CP-element group 359:  members (12) 
      -- CP-element group 359: 	 branch_block_stmt_26/if_stmt_1279_else_link/$exit
      -- CP-element group 359: 	 branch_block_stmt_26/if_stmt_1279_else_link/else_choice_transition
      -- CP-element group 359: 	 branch_block_stmt_26/forx_xbody370_forx_xbody370
      -- CP-element group 359: 	 branch_block_stmt_26/forx_xbody370_forx_xbody370_PhiReq/$entry
      -- CP-element group 359: 	 branch_block_stmt_26/forx_xbody370_forx_xbody370_PhiReq/phi_stmt_1151/$entry
      -- CP-element group 359: 	 branch_block_stmt_26/forx_xbody370_forx_xbody370_PhiReq/phi_stmt_1151/phi_stmt_1151_sources/$entry
      -- CP-element group 359: 	 branch_block_stmt_26/forx_xbody370_forx_xbody370_PhiReq/phi_stmt_1151/phi_stmt_1151_sources/type_cast_1157/$entry
      -- CP-element group 359: 	 branch_block_stmt_26/forx_xbody370_forx_xbody370_PhiReq/phi_stmt_1151/phi_stmt_1151_sources/type_cast_1157/SplitProtocol/$entry
      -- CP-element group 359: 	 branch_block_stmt_26/forx_xbody370_forx_xbody370_PhiReq/phi_stmt_1151/phi_stmt_1151_sources/type_cast_1157/SplitProtocol/Sample/$entry
      -- CP-element group 359: 	 branch_block_stmt_26/forx_xbody370_forx_xbody370_PhiReq/phi_stmt_1151/phi_stmt_1151_sources/type_cast_1157/SplitProtocol/Sample/rr
      -- CP-element group 359: 	 branch_block_stmt_26/forx_xbody370_forx_xbody370_PhiReq/phi_stmt_1151/phi_stmt_1151_sources/type_cast_1157/SplitProtocol/Update/$entry
      -- CP-element group 359: 	 branch_block_stmt_26/forx_xbody370_forx_xbody370_PhiReq/phi_stmt_1151/phi_stmt_1151_sources/type_cast_1157/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 359_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1279_branch_ack_0, ack => convTranspose_CP_39_elements(359)); -- 
    rr_3010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(359), ack => type_cast_1157_inst_req_0); -- 
    cr_3015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(359), ack => type_cast_1157_inst_req_1); -- 
    -- CP-element group 360:  merge  branch  transition  place  output  bypass 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	165 
    -- CP-element group 360: 	120 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	121 
    -- CP-element group 360: 	122 
    -- CP-element group 360:  members (17) 
      -- CP-element group 360: 	 branch_block_stmt_26/merge_stmt_395__exit__
      -- CP-element group 360: 	 branch_block_stmt_26/assign_stmt_401__entry__
      -- CP-element group 360: 	 branch_block_stmt_26/assign_stmt_401__exit__
      -- CP-element group 360: 	 branch_block_stmt_26/if_stmt_402__entry__
      -- CP-element group 360: 	 branch_block_stmt_26/assign_stmt_401/$entry
      -- CP-element group 360: 	 branch_block_stmt_26/assign_stmt_401/$exit
      -- CP-element group 360: 	 branch_block_stmt_26/if_stmt_402_dead_link/$entry
      -- CP-element group 360: 	 branch_block_stmt_26/if_stmt_402_eval_test/$entry
      -- CP-element group 360: 	 branch_block_stmt_26/if_stmt_402_eval_test/$exit
      -- CP-element group 360: 	 branch_block_stmt_26/if_stmt_402_eval_test/branch_req
      -- CP-element group 360: 	 branch_block_stmt_26/R_cmp194452_403_place
      -- CP-element group 360: 	 branch_block_stmt_26/if_stmt_402_if_link/$entry
      -- CP-element group 360: 	 branch_block_stmt_26/if_stmt_402_else_link/$entry
      -- CP-element group 360: 	 branch_block_stmt_26/merge_stmt_395_PhiReqMerge
      -- CP-element group 360: 	 branch_block_stmt_26/merge_stmt_395_PhiAck/$entry
      -- CP-element group 360: 	 branch_block_stmt_26/merge_stmt_395_PhiAck/$exit
      -- CP-element group 360: 	 branch_block_stmt_26/merge_stmt_395_PhiAck/dummy
      -- 
    branch_req_929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(360), ack => if_stmt_402_branch_req_0); -- 
    convTranspose_CP_39_elements(360) <= OrReduce(convTranspose_CP_39_elements(165) & convTranspose_CP_39_elements(120));
    -- CP-element group 361:  transition  output  delay-element  bypass 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	124 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	365 
    -- CP-element group 361:  members (5) 
      -- CP-element group 361: 	 branch_block_stmt_26/bbx_xnph458_forx_xbody_PhiReq/$exit
      -- CP-element group 361: 	 branch_block_stmt_26/bbx_xnph458_forx_xbody_PhiReq/phi_stmt_446/$exit
      -- CP-element group 361: 	 branch_block_stmt_26/bbx_xnph458_forx_xbody_PhiReq/phi_stmt_446/phi_stmt_446_sources/$exit
      -- CP-element group 361: 	 branch_block_stmt_26/bbx_xnph458_forx_xbody_PhiReq/phi_stmt_446/phi_stmt_446_sources/type_cast_450_konst_delay_trans
      -- CP-element group 361: 	 branch_block_stmt_26/bbx_xnph458_forx_xbody_PhiReq/phi_stmt_446/phi_stmt_446_req
      -- 
    phi_stmt_446_req_2783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_446_req_2783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(361), ack => phi_stmt_446_req_0); -- 
    -- Element group convTranspose_CP_39_elements(361) is a control-delay.
    cp_element_361_delay: control_delay_element  generic map(name => " 361_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(124), ack => convTranspose_CP_39_elements(361), clk => clk, reset =>reset);
    -- CP-element group 362:  transition  input  bypass 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	166 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	364 
    -- CP-element group 362:  members (2) 
      -- CP-element group 362: 	 branch_block_stmt_26/forx_xbody_forx_xbody_PhiReq/phi_stmt_446/phi_stmt_446_sources/type_cast_452/SplitProtocol/Sample/$exit
      -- CP-element group 362: 	 branch_block_stmt_26/forx_xbody_forx_xbody_PhiReq/phi_stmt_446/phi_stmt_446_sources/type_cast_452/SplitProtocol/Sample/ra
      -- 
    ra_2803_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 362_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_452_inst_ack_0, ack => convTranspose_CP_39_elements(362)); -- 
    -- CP-element group 363:  transition  input  bypass 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	166 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	364 
    -- CP-element group 363:  members (2) 
      -- CP-element group 363: 	 branch_block_stmt_26/forx_xbody_forx_xbody_PhiReq/phi_stmt_446/phi_stmt_446_sources/type_cast_452/SplitProtocol/Update/$exit
      -- CP-element group 363: 	 branch_block_stmt_26/forx_xbody_forx_xbody_PhiReq/phi_stmt_446/phi_stmt_446_sources/type_cast_452/SplitProtocol/Update/ca
      -- 
    ca_2808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 363_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_452_inst_ack_1, ack => convTranspose_CP_39_elements(363)); -- 
    -- CP-element group 364:  join  transition  output  bypass 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	362 
    -- CP-element group 364: 	363 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	365 
    -- CP-element group 364:  members (6) 
      -- CP-element group 364: 	 branch_block_stmt_26/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 364: 	 branch_block_stmt_26/forx_xbody_forx_xbody_PhiReq/phi_stmt_446/$exit
      -- CP-element group 364: 	 branch_block_stmt_26/forx_xbody_forx_xbody_PhiReq/phi_stmt_446/phi_stmt_446_sources/$exit
      -- CP-element group 364: 	 branch_block_stmt_26/forx_xbody_forx_xbody_PhiReq/phi_stmt_446/phi_stmt_446_sources/type_cast_452/$exit
      -- CP-element group 364: 	 branch_block_stmt_26/forx_xbody_forx_xbody_PhiReq/phi_stmt_446/phi_stmt_446_sources/type_cast_452/SplitProtocol/$exit
      -- CP-element group 364: 	 branch_block_stmt_26/forx_xbody_forx_xbody_PhiReq/phi_stmt_446/phi_stmt_446_req
      -- 
    phi_stmt_446_req_2809_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_446_req_2809_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(364), ack => phi_stmt_446_req_1); -- 
    convTranspose_cp_element_group_364: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_364"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(362) & convTranspose_CP_39_elements(363);
      gj_convTranspose_cp_element_group_364 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(364), clk => clk, reset => reset); --
    end block;
    -- CP-element group 365:  merge  transition  place  bypass 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	361 
    -- CP-element group 365: 	364 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	366 
    -- CP-element group 365:  members (2) 
      -- CP-element group 365: 	 branch_block_stmt_26/merge_stmt_445_PhiReqMerge
      -- CP-element group 365: 	 branch_block_stmt_26/merge_stmt_445_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(365) <= OrReduce(convTranspose_CP_39_elements(361) & convTranspose_CP_39_elements(364));
    -- CP-element group 366:  fork  transition  place  input  output  bypass 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	365 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	136 
    -- CP-element group 366: 	140 
    -- CP-element group 366: 	129 
    -- CP-element group 366: 	132 
    -- CP-element group 366: 	144 
    -- CP-element group 366: 	148 
    -- CP-element group 366: 	152 
    -- CP-element group 366: 	156 
    -- CP-element group 366: 	160 
    -- CP-element group 366: 	163 
    -- CP-element group 366: 	125 
    -- CP-element group 366: 	126 
    -- CP-element group 366: 	128 
    -- CP-element group 366:  members (56) 
      -- CP-element group 366: 	 branch_block_stmt_26/merge_stmt_445__exit__
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608__entry__
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_569_Update/cr
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_569_Update/$entry
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_515_Update/cr
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_515_Update/$entry
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/ptr_deref_595_Update/$entry
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/ptr_deref_595_update_start_
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/ptr_deref_595_Update/word_access_complete/word_0/cr
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/ptr_deref_595_Update/word_access_complete/word_0/$entry
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/ptr_deref_595_Update/word_access_complete/$entry
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_569_update_start_
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_551_Update/cr
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_551_Update/$entry
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_587_Update/cr
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_587_Update/$entry
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_515_update_start_
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_551_update_start_
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_587_update_start_
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_533_Update/cr
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_533_Update/$entry
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_533_update_start_
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/$entry
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/addr_of_459_update_start_
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/array_obj_ref_458_index_resized_1
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/array_obj_ref_458_index_scaled_1
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/array_obj_ref_458_index_computed_1
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/array_obj_ref_458_index_resize_1/$entry
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/array_obj_ref_458_index_resize_1/$exit
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/array_obj_ref_458_index_resize_1/index_resize_req
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/array_obj_ref_458_index_resize_1/index_resize_ack
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/array_obj_ref_458_index_scale_1/$entry
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/array_obj_ref_458_index_scale_1/$exit
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/array_obj_ref_458_index_scale_1/scale_rename_req
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/array_obj_ref_458_index_scale_1/scale_rename_ack
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/array_obj_ref_458_final_index_sum_regn_update_start
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/array_obj_ref_458_final_index_sum_regn_Sample/$entry
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/array_obj_ref_458_final_index_sum_regn_Sample/req
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/array_obj_ref_458_final_index_sum_regn_Update/$entry
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/array_obj_ref_458_final_index_sum_regn_Update/req
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/addr_of_459_complete/$entry
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/addr_of_459_complete/req
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_462_sample_start_
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_462_Sample/$entry
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/RPIPE_ConvTranspose_input_pipe_462_Sample/rr
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_466_update_start_
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_466_Update/$entry
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_466_Update/cr
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_479_update_start_
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_479_Update/$entry
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_479_Update/cr
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_497_update_start_
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_497_Update/$entry
      -- CP-element group 366: 	 branch_block_stmt_26/assign_stmt_460_to_assign_stmt_608/type_cast_497_Update/cr
      -- CP-element group 366: 	 branch_block_stmt_26/merge_stmt_445_PhiAck/$exit
      -- CP-element group 366: 	 branch_block_stmt_26/merge_stmt_445_PhiAck/phi_stmt_446_ack
      -- 
    phi_stmt_446_ack_2814_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 366_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_446_ack_0, ack => convTranspose_CP_39_elements(366)); -- 
    cr_1201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(366), ack => type_cast_569_inst_req_1); -- 
    cr_1117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(366), ack => type_cast_515_inst_req_1); -- 
    cr_1279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(366), ack => ptr_deref_595_store_0_req_1); -- 
    cr_1173_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1173_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(366), ack => type_cast_551_inst_req_1); -- 
    cr_1229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(366), ack => type_cast_587_inst_req_1); -- 
    cr_1145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(366), ack => type_cast_533_inst_req_1); -- 
    req_985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(366), ack => array_obj_ref_458_index_offset_req_0); -- 
    req_990_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_990_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(366), ack => array_obj_ref_458_index_offset_req_1); -- 
    req_1005_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1005_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(366), ack => addr_of_459_final_reg_req_1); -- 
    rr_1014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(366), ack => RPIPE_ConvTranspose_input_pipe_462_inst_req_0); -- 
    cr_1033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(366), ack => type_cast_466_inst_req_1); -- 
    cr_1061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(366), ack => type_cast_479_inst_req_1); -- 
    cr_1089_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1089_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(366), ack => type_cast_497_inst_req_1); -- 
    -- CP-element group 367:  transition  output  delay-element  bypass 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	168 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	371 
    -- CP-element group 367:  members (5) 
      -- CP-element group 367: 	 branch_block_stmt_26/bbx_xnph454_forx_xbody196_PhiReq/$exit
      -- CP-element group 367: 	 branch_block_stmt_26/bbx_xnph454_forx_xbody196_PhiReq/phi_stmt_653/$exit
      -- CP-element group 367: 	 branch_block_stmt_26/bbx_xnph454_forx_xbody196_PhiReq/phi_stmt_653/phi_stmt_653_sources/$exit
      -- CP-element group 367: 	 branch_block_stmt_26/bbx_xnph454_forx_xbody196_PhiReq/phi_stmt_653/phi_stmt_653_sources/type_cast_657_konst_delay_trans
      -- CP-element group 367: 	 branch_block_stmt_26/bbx_xnph454_forx_xbody196_PhiReq/phi_stmt_653/phi_stmt_653_req
      -- 
    phi_stmt_653_req_2837_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_653_req_2837_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(367), ack => phi_stmt_653_req_0); -- 
    -- Element group convTranspose_CP_39_elements(367) is a control-delay.
    cp_element_367_delay: control_delay_element  generic map(name => " 367_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(168), ack => convTranspose_CP_39_elements(367), clk => clk, reset =>reset);
    -- CP-element group 368:  transition  input  bypass 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	210 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	370 
    -- CP-element group 368:  members (2) 
      -- CP-element group 368: 	 branch_block_stmt_26/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_653/phi_stmt_653_sources/type_cast_659/SplitProtocol/Sample/$exit
      -- CP-element group 368: 	 branch_block_stmt_26/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_653/phi_stmt_653_sources/type_cast_659/SplitProtocol/Sample/ra
      -- 
    ra_2857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 368_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_659_inst_ack_0, ack => convTranspose_CP_39_elements(368)); -- 
    -- CP-element group 369:  transition  input  bypass 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	210 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	370 
    -- CP-element group 369:  members (2) 
      -- CP-element group 369: 	 branch_block_stmt_26/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_653/phi_stmt_653_sources/type_cast_659/SplitProtocol/Update/$exit
      -- CP-element group 369: 	 branch_block_stmt_26/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_653/phi_stmt_653_sources/type_cast_659/SplitProtocol/Update/ca
      -- 
    ca_2862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 369_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_659_inst_ack_1, ack => convTranspose_CP_39_elements(369)); -- 
    -- CP-element group 370:  join  transition  output  bypass 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	368 
    -- CP-element group 370: 	369 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	371 
    -- CP-element group 370:  members (6) 
      -- CP-element group 370: 	 branch_block_stmt_26/forx_xbody196_forx_xbody196_PhiReq/$exit
      -- CP-element group 370: 	 branch_block_stmt_26/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_653/$exit
      -- CP-element group 370: 	 branch_block_stmt_26/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_653/phi_stmt_653_sources/$exit
      -- CP-element group 370: 	 branch_block_stmt_26/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_653/phi_stmt_653_sources/type_cast_659/$exit
      -- CP-element group 370: 	 branch_block_stmt_26/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_653/phi_stmt_653_sources/type_cast_659/SplitProtocol/$exit
      -- CP-element group 370: 	 branch_block_stmt_26/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_653/phi_stmt_653_req
      -- 
    phi_stmt_653_req_2863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_653_req_2863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(370), ack => phi_stmt_653_req_1); -- 
    convTranspose_cp_element_group_370: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_370"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(368) & convTranspose_CP_39_elements(369);
      gj_convTranspose_cp_element_group_370 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(370), clk => clk, reset => reset); --
    end block;
    -- CP-element group 371:  merge  transition  place  bypass 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	367 
    -- CP-element group 371: 	370 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	372 
    -- CP-element group 371:  members (2) 
      -- CP-element group 371: 	 branch_block_stmt_26/merge_stmt_652_PhiReqMerge
      -- CP-element group 371: 	 branch_block_stmt_26/merge_stmt_652_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(371) <= OrReduce(convTranspose_CP_39_elements(367) & convTranspose_CP_39_elements(370));
    -- CP-element group 372:  fork  transition  place  input  output  bypass 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	371 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	169 
    -- CP-element group 372: 	170 
    -- CP-element group 372: 	172 
    -- CP-element group 372: 	173 
    -- CP-element group 372: 	176 
    -- CP-element group 372: 	180 
    -- CP-element group 372: 	184 
    -- CP-element group 372: 	188 
    -- CP-element group 372: 	192 
    -- CP-element group 372: 	196 
    -- CP-element group 372: 	200 
    -- CP-element group 372: 	204 
    -- CP-element group 372: 	207 
    -- CP-element group 372:  members (56) 
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_722_update_start_
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/array_obj_ref_665_index_resize_1/$entry
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_704_update_start_
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/array_obj_ref_665_index_resize_1/$exit
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_669_sample_start_
      -- CP-element group 372: 	 branch_block_stmt_26/merge_stmt_652__exit__
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815__entry__
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_686_update_start_
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_686_Update/cr
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_673_update_start_
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/array_obj_ref_665_index_resize_1/index_resize_ack
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/array_obj_ref_665_index_computed_1
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_704_Update/cr
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/addr_of_666_update_start_
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_686_Update/$entry
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/array_obj_ref_665_index_scaled_1
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_704_Update/$entry
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/$entry
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/array_obj_ref_665_index_resized_1
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_669_Sample/rr
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/RPIPE_ConvTranspose_input_pipe_669_Sample/$entry
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/array_obj_ref_665_index_resize_1/index_resize_req
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/array_obj_ref_665_final_index_sum_regn_Update/req
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/array_obj_ref_665_final_index_sum_regn_Update/$entry
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/array_obj_ref_665_final_index_sum_regn_Sample/req
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/array_obj_ref_665_final_index_sum_regn_Sample/$entry
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/array_obj_ref_665_final_index_sum_regn_update_start
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/array_obj_ref_665_index_scale_1/scale_rename_ack
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/array_obj_ref_665_index_scale_1/scale_rename_req
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_673_Update/cr
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/addr_of_666_complete/req
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/array_obj_ref_665_index_scale_1/$exit
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/array_obj_ref_665_index_scale_1/$entry
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_673_Update/$entry
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/addr_of_666_complete/$entry
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_722_Update/$entry
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_722_Update/cr
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_740_update_start_
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_740_Update/$entry
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_740_Update/cr
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_758_update_start_
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_758_Update/$entry
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_758_Update/cr
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_776_update_start_
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_776_Update/$entry
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_776_Update/cr
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_794_update_start_
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_794_Update/$entry
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/type_cast_794_Update/cr
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/ptr_deref_802_update_start_
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/ptr_deref_802_Update/$entry
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/ptr_deref_802_Update/word_access_complete/$entry
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/ptr_deref_802_Update/word_access_complete/word_0/$entry
      -- CP-element group 372: 	 branch_block_stmt_26/assign_stmt_667_to_assign_stmt_815/ptr_deref_802_Update/word_access_complete/word_0/cr
      -- CP-element group 372: 	 branch_block_stmt_26/merge_stmt_652_PhiAck/$exit
      -- CP-element group 372: 	 branch_block_stmt_26/merge_stmt_652_PhiAck/phi_stmt_653_ack
      -- 
    phi_stmt_653_ack_2868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 372_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_653_ack_0, ack => convTranspose_CP_39_elements(372)); -- 
    cr_1420_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1420_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(372), ack => type_cast_686_inst_req_1); -- 
    cr_1448_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1448_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(372), ack => type_cast_704_inst_req_1); -- 
    rr_1373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(372), ack => RPIPE_ConvTranspose_input_pipe_669_inst_req_0); -- 
    req_1349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(372), ack => array_obj_ref_665_index_offset_req_1); -- 
    req_1344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(372), ack => array_obj_ref_665_index_offset_req_0); -- 
    cr_1392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(372), ack => type_cast_673_inst_req_1); -- 
    req_1364_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1364_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(372), ack => addr_of_666_final_reg_req_1); -- 
    cr_1476_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1476_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(372), ack => type_cast_722_inst_req_1); -- 
    cr_1504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(372), ack => type_cast_740_inst_req_1); -- 
    cr_1532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(372), ack => type_cast_758_inst_req_1); -- 
    cr_1560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(372), ack => type_cast_776_inst_req_1); -- 
    cr_1588_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1588_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(372), ack => type_cast_794_inst_req_1); -- 
    cr_1638_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1638_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(372), ack => ptr_deref_802_store_0_req_1); -- 
    -- CP-element group 373:  merge  fork  transition  place  output  bypass 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	209 
    -- CP-element group 373: 	122 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	211 
    -- CP-element group 373: 	212 
    -- CP-element group 373: 	213 
    -- CP-element group 373: 	214 
    -- CP-element group 373: 	215 
    -- CP-element group 373: 	216 
    -- CP-element group 373:  members (25) 
      -- CP-element group 373: 	 branch_block_stmt_26/merge_stmt_824__exit__
      -- CP-element group 373: 	 branch_block_stmt_26/assign_stmt_828_to_assign_stmt_852__entry__
      -- CP-element group 373: 	 branch_block_stmt_26/assign_stmt_828_to_assign_stmt_852/$entry
      -- CP-element group 373: 	 branch_block_stmt_26/assign_stmt_828_to_assign_stmt_852/type_cast_827_sample_start_
      -- CP-element group 373: 	 branch_block_stmt_26/assign_stmt_828_to_assign_stmt_852/type_cast_827_update_start_
      -- CP-element group 373: 	 branch_block_stmt_26/assign_stmt_828_to_assign_stmt_852/type_cast_827_Sample/$entry
      -- CP-element group 373: 	 branch_block_stmt_26/assign_stmt_828_to_assign_stmt_852/type_cast_827_Sample/rr
      -- CP-element group 373: 	 branch_block_stmt_26/assign_stmt_828_to_assign_stmt_852/type_cast_827_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_26/assign_stmt_828_to_assign_stmt_852/type_cast_827_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_26/assign_stmt_828_to_assign_stmt_852/type_cast_831_sample_start_
      -- CP-element group 373: 	 branch_block_stmt_26/assign_stmt_828_to_assign_stmt_852/type_cast_831_update_start_
      -- CP-element group 373: 	 branch_block_stmt_26/assign_stmt_828_to_assign_stmt_852/type_cast_831_Sample/$entry
      -- CP-element group 373: 	 branch_block_stmt_26/assign_stmt_828_to_assign_stmt_852/type_cast_831_Sample/rr
      -- CP-element group 373: 	 branch_block_stmt_26/assign_stmt_828_to_assign_stmt_852/type_cast_831_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_26/assign_stmt_828_to_assign_stmt_852/type_cast_831_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_26/assign_stmt_828_to_assign_stmt_852/type_cast_835_sample_start_
      -- CP-element group 373: 	 branch_block_stmt_26/assign_stmt_828_to_assign_stmt_852/type_cast_835_update_start_
      -- CP-element group 373: 	 branch_block_stmt_26/assign_stmt_828_to_assign_stmt_852/type_cast_835_Sample/$entry
      -- CP-element group 373: 	 branch_block_stmt_26/assign_stmt_828_to_assign_stmt_852/type_cast_835_Sample/rr
      -- CP-element group 373: 	 branch_block_stmt_26/assign_stmt_828_to_assign_stmt_852/type_cast_835_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_26/assign_stmt_828_to_assign_stmt_852/type_cast_835_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_26/merge_stmt_824_PhiReqMerge
      -- CP-element group 373: 	 branch_block_stmt_26/merge_stmt_824_PhiAck/$entry
      -- CP-element group 373: 	 branch_block_stmt_26/merge_stmt_824_PhiAck/$exit
      -- CP-element group 373: 	 branch_block_stmt_26/merge_stmt_824_PhiAck/dummy
      -- 
    rr_1669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => type_cast_827_inst_req_0); -- 
    cr_1674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => type_cast_827_inst_req_1); -- 
    rr_1683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => type_cast_831_inst_req_0); -- 
    cr_1688_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1688_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => type_cast_831_inst_req_1); -- 
    rr_1697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => type_cast_835_inst_req_0); -- 
    cr_1702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => type_cast_835_inst_req_1); -- 
    convTranspose_CP_39_elements(373) <= OrReduce(convTranspose_CP_39_elements(209) & convTranspose_CP_39_elements(122));
    -- CP-element group 374:  transition  output  delay-element  bypass 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	221 
    -- CP-element group 374: successors 
    -- CP-element group 374: 	378 
    -- CP-element group 374:  members (5) 
      -- CP-element group 374: 	 branch_block_stmt_26/bbx_xnph450_forx_xbody266_PhiReq/$exit
      -- CP-element group 374: 	 branch_block_stmt_26/bbx_xnph450_forx_xbody266_PhiReq/phi_stmt_897/$exit
      -- CP-element group 374: 	 branch_block_stmt_26/bbx_xnph450_forx_xbody266_PhiReq/phi_stmt_897/phi_stmt_897_sources/$exit
      -- CP-element group 374: 	 branch_block_stmt_26/bbx_xnph450_forx_xbody266_PhiReq/phi_stmt_897/phi_stmt_897_sources/type_cast_901_konst_delay_trans
      -- CP-element group 374: 	 branch_block_stmt_26/bbx_xnph450_forx_xbody266_PhiReq/phi_stmt_897/phi_stmt_897_req
      -- 
    phi_stmt_897_req_2914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_897_req_2914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(374), ack => phi_stmt_897_req_0); -- 
    -- Element group convTranspose_CP_39_elements(374) is a control-delay.
    cp_element_374_delay: control_delay_element  generic map(name => " 374_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(221), ack => convTranspose_CP_39_elements(374), clk => clk, reset =>reset);
    -- CP-element group 375:  transition  input  bypass 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	230 
    -- CP-element group 375: successors 
    -- CP-element group 375: 	377 
    -- CP-element group 375:  members (2) 
      -- CP-element group 375: 	 branch_block_stmt_26/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_897/phi_stmt_897_sources/type_cast_903/SplitProtocol/Sample/$exit
      -- CP-element group 375: 	 branch_block_stmt_26/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_897/phi_stmt_897_sources/type_cast_903/SplitProtocol/Sample/ra
      -- 
    ra_2934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 375_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_903_inst_ack_0, ack => convTranspose_CP_39_elements(375)); -- 
    -- CP-element group 376:  transition  input  bypass 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	230 
    -- CP-element group 376: successors 
    -- CP-element group 376: 	377 
    -- CP-element group 376:  members (2) 
      -- CP-element group 376: 	 branch_block_stmt_26/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_897/phi_stmt_897_sources/type_cast_903/SplitProtocol/Update/$exit
      -- CP-element group 376: 	 branch_block_stmt_26/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_897/phi_stmt_897_sources/type_cast_903/SplitProtocol/Update/ca
      -- 
    ca_2939_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 376_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_903_inst_ack_1, ack => convTranspose_CP_39_elements(376)); -- 
    -- CP-element group 377:  join  transition  output  bypass 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	375 
    -- CP-element group 377: 	376 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	378 
    -- CP-element group 377:  members (6) 
      -- CP-element group 377: 	 branch_block_stmt_26/forx_xbody266_forx_xbody266_PhiReq/$exit
      -- CP-element group 377: 	 branch_block_stmt_26/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_897/$exit
      -- CP-element group 377: 	 branch_block_stmt_26/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_897/phi_stmt_897_sources/$exit
      -- CP-element group 377: 	 branch_block_stmt_26/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_897/phi_stmt_897_sources/type_cast_903/$exit
      -- CP-element group 377: 	 branch_block_stmt_26/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_897/phi_stmt_897_sources/type_cast_903/SplitProtocol/$exit
      -- CP-element group 377: 	 branch_block_stmt_26/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_897/phi_stmt_897_req
      -- 
    phi_stmt_897_req_2940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_897_req_2940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(377), ack => phi_stmt_897_req_1); -- 
    convTranspose_cp_element_group_377: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_377"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(375) & convTranspose_CP_39_elements(376);
      gj_convTranspose_cp_element_group_377 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(377), clk => clk, reset => reset); --
    end block;
    -- CP-element group 378:  merge  transition  place  bypass 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	374 
    -- CP-element group 378: 	377 
    -- CP-element group 378: successors 
    -- CP-element group 378: 	379 
    -- CP-element group 378:  members (2) 
      -- CP-element group 378: 	 branch_block_stmt_26/merge_stmt_896_PhiReqMerge
      -- CP-element group 378: 	 branch_block_stmt_26/merge_stmt_896_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(378) <= OrReduce(convTranspose_CP_39_elements(374) & convTranspose_CP_39_elements(377));
    -- CP-element group 379:  fork  transition  place  input  output  bypass 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	378 
    -- CP-element group 379: successors 
    -- CP-element group 379: 	222 
    -- CP-element group 379: 	223 
    -- CP-element group 379: 	225 
    -- CP-element group 379: 	227 
    -- CP-element group 379:  members (29) 
      -- CP-element group 379: 	 branch_block_stmt_26/merge_stmt_896__exit__
      -- CP-element group 379: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927__entry__
      -- CP-element group 379: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/$entry
      -- CP-element group 379: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/addr_of_910_update_start_
      -- CP-element group 379: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/array_obj_ref_909_index_resized_1
      -- CP-element group 379: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/array_obj_ref_909_index_scaled_1
      -- CP-element group 379: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/array_obj_ref_909_index_computed_1
      -- CP-element group 379: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/array_obj_ref_909_index_resize_1/$entry
      -- CP-element group 379: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/array_obj_ref_909_index_resize_1/$exit
      -- CP-element group 379: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/array_obj_ref_909_index_resize_1/index_resize_req
      -- CP-element group 379: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/array_obj_ref_909_index_resize_1/index_resize_ack
      -- CP-element group 379: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/array_obj_ref_909_index_scale_1/$entry
      -- CP-element group 379: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/array_obj_ref_909_index_scale_1/$exit
      -- CP-element group 379: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/array_obj_ref_909_index_scale_1/scale_rename_req
      -- CP-element group 379: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/array_obj_ref_909_index_scale_1/scale_rename_ack
      -- CP-element group 379: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/array_obj_ref_909_final_index_sum_regn_update_start
      -- CP-element group 379: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/array_obj_ref_909_final_index_sum_regn_Sample/$entry
      -- CP-element group 379: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/array_obj_ref_909_final_index_sum_regn_Sample/req
      -- CP-element group 379: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/array_obj_ref_909_final_index_sum_regn_Update/$entry
      -- CP-element group 379: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/array_obj_ref_909_final_index_sum_regn_Update/req
      -- CP-element group 379: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/addr_of_910_complete/$entry
      -- CP-element group 379: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/addr_of_910_complete/req
      -- CP-element group 379: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/ptr_deref_913_update_start_
      -- CP-element group 379: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/ptr_deref_913_Update/$entry
      -- CP-element group 379: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/ptr_deref_913_Update/word_access_complete/$entry
      -- CP-element group 379: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/ptr_deref_913_Update/word_access_complete/word_0/$entry
      -- CP-element group 379: 	 branch_block_stmt_26/assign_stmt_911_to_assign_stmt_927/ptr_deref_913_Update/word_access_complete/word_0/cr
      -- CP-element group 379: 	 branch_block_stmt_26/merge_stmt_896_PhiAck/$exit
      -- CP-element group 379: 	 branch_block_stmt_26/merge_stmt_896_PhiAck/phi_stmt_897_ack
      -- 
    phi_stmt_897_ack_2945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 379_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_897_ack_0, ack => convTranspose_CP_39_elements(379)); -- 
    req_1767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(379), ack => array_obj_ref_909_index_offset_req_0); -- 
    req_1772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(379), ack => array_obj_ref_909_index_offset_req_1); -- 
    req_1787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(379), ack => addr_of_910_final_reg_req_1); -- 
    cr_1837_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1837_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(379), ack => ptr_deref_913_store_0_req_1); -- 
    -- CP-element group 380:  merge  fork  transition  place  output  bypass 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	219 
    -- CP-element group 380: 	229 
    -- CP-element group 380: successors 
    -- CP-element group 380: 	231 
    -- CP-element group 380: 	232 
    -- CP-element group 380: 	234 
    -- CP-element group 380:  members (16) 
      -- CP-element group 380: 	 branch_block_stmt_26/merge_stmt_936__exit__
      -- CP-element group 380: 	 branch_block_stmt_26/call_stmt_939_to_assign_stmt_945__entry__
      -- CP-element group 380: 	 branch_block_stmt_26/call_stmt_939_to_assign_stmt_945/$entry
      -- CP-element group 380: 	 branch_block_stmt_26/call_stmt_939_to_assign_stmt_945/call_stmt_939_sample_start_
      -- CP-element group 380: 	 branch_block_stmt_26/call_stmt_939_to_assign_stmt_945/call_stmt_939_update_start_
      -- CP-element group 380: 	 branch_block_stmt_26/call_stmt_939_to_assign_stmt_945/call_stmt_939_Sample/$entry
      -- CP-element group 380: 	 branch_block_stmt_26/call_stmt_939_to_assign_stmt_945/call_stmt_939_Sample/crr
      -- CP-element group 380: 	 branch_block_stmt_26/call_stmt_939_to_assign_stmt_945/call_stmt_939_Update/$entry
      -- CP-element group 380: 	 branch_block_stmt_26/call_stmt_939_to_assign_stmt_945/call_stmt_939_Update/ccr
      -- CP-element group 380: 	 branch_block_stmt_26/call_stmt_939_to_assign_stmt_945/type_cast_944_update_start_
      -- CP-element group 380: 	 branch_block_stmt_26/call_stmt_939_to_assign_stmt_945/type_cast_944_Update/$entry
      -- CP-element group 380: 	 branch_block_stmt_26/call_stmt_939_to_assign_stmt_945/type_cast_944_Update/cr
      -- CP-element group 380: 	 branch_block_stmt_26/merge_stmt_936_PhiReqMerge
      -- CP-element group 380: 	 branch_block_stmt_26/merge_stmt_936_PhiAck/$entry
      -- CP-element group 380: 	 branch_block_stmt_26/merge_stmt_936_PhiAck/$exit
      -- CP-element group 380: 	 branch_block_stmt_26/merge_stmt_936_PhiAck/dummy
      -- 
    crr_1868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(380), ack => call_stmt_939_call_req_0); -- 
    ccr_1873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(380), ack => call_stmt_939_call_req_1); -- 
    cr_1887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(380), ack => type_cast_944_inst_req_1); -- 
    convTranspose_CP_39_elements(380) <= OrReduce(convTranspose_CP_39_elements(219) & convTranspose_CP_39_elements(229));
    -- CP-element group 381:  transition  output  delay-element  bypass 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	311 
    -- CP-element group 381: successors 
    -- CP-element group 381: 	385 
    -- CP-element group 381:  members (5) 
      -- CP-element group 381: 	 branch_block_stmt_26/bbx_xnph_forx_xbody370_PhiReq/$exit
      -- CP-element group 381: 	 branch_block_stmt_26/bbx_xnph_forx_xbody370_PhiReq/phi_stmt_1151/$exit
      -- CP-element group 381: 	 branch_block_stmt_26/bbx_xnph_forx_xbody370_PhiReq/phi_stmt_1151/phi_stmt_1151_sources/$exit
      -- CP-element group 381: 	 branch_block_stmt_26/bbx_xnph_forx_xbody370_PhiReq/phi_stmt_1151/phi_stmt_1151_sources/type_cast_1155_konst_delay_trans
      -- CP-element group 381: 	 branch_block_stmt_26/bbx_xnph_forx_xbody370_PhiReq/phi_stmt_1151/phi_stmt_1151_req
      -- 
    phi_stmt_1151_req_2991_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1151_req_2991_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(381), ack => phi_stmt_1151_req_0); -- 
    -- Element group convTranspose_CP_39_elements(381) is a control-delay.
    cp_element_381_delay: control_delay_element  generic map(name => " 381_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(311), ack => convTranspose_CP_39_elements(381), clk => clk, reset =>reset);
    -- CP-element group 382:  transition  input  bypass 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	359 
    -- CP-element group 382: successors 
    -- CP-element group 382: 	384 
    -- CP-element group 382:  members (2) 
      -- CP-element group 382: 	 branch_block_stmt_26/forx_xbody370_forx_xbody370_PhiReq/phi_stmt_1151/phi_stmt_1151_sources/type_cast_1157/SplitProtocol/Sample/$exit
      -- CP-element group 382: 	 branch_block_stmt_26/forx_xbody370_forx_xbody370_PhiReq/phi_stmt_1151/phi_stmt_1151_sources/type_cast_1157/SplitProtocol/Sample/ra
      -- 
    ra_3011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 382_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1157_inst_ack_0, ack => convTranspose_CP_39_elements(382)); -- 
    -- CP-element group 383:  transition  input  bypass 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	359 
    -- CP-element group 383: successors 
    -- CP-element group 383: 	384 
    -- CP-element group 383:  members (2) 
      -- CP-element group 383: 	 branch_block_stmt_26/forx_xbody370_forx_xbody370_PhiReq/phi_stmt_1151/phi_stmt_1151_sources/type_cast_1157/SplitProtocol/Update/$exit
      -- CP-element group 383: 	 branch_block_stmt_26/forx_xbody370_forx_xbody370_PhiReq/phi_stmt_1151/phi_stmt_1151_sources/type_cast_1157/SplitProtocol/Update/ca
      -- 
    ca_3016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 383_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1157_inst_ack_1, ack => convTranspose_CP_39_elements(383)); -- 
    -- CP-element group 384:  join  transition  output  bypass 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	382 
    -- CP-element group 384: 	383 
    -- CP-element group 384: successors 
    -- CP-element group 384: 	385 
    -- CP-element group 384:  members (6) 
      -- CP-element group 384: 	 branch_block_stmt_26/forx_xbody370_forx_xbody370_PhiReq/$exit
      -- CP-element group 384: 	 branch_block_stmt_26/forx_xbody370_forx_xbody370_PhiReq/phi_stmt_1151/$exit
      -- CP-element group 384: 	 branch_block_stmt_26/forx_xbody370_forx_xbody370_PhiReq/phi_stmt_1151/phi_stmt_1151_sources/$exit
      -- CP-element group 384: 	 branch_block_stmt_26/forx_xbody370_forx_xbody370_PhiReq/phi_stmt_1151/phi_stmt_1151_sources/type_cast_1157/$exit
      -- CP-element group 384: 	 branch_block_stmt_26/forx_xbody370_forx_xbody370_PhiReq/phi_stmt_1151/phi_stmt_1151_sources/type_cast_1157/SplitProtocol/$exit
      -- CP-element group 384: 	 branch_block_stmt_26/forx_xbody370_forx_xbody370_PhiReq/phi_stmt_1151/phi_stmt_1151_req
      -- 
    phi_stmt_1151_req_3017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1151_req_3017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(384), ack => phi_stmt_1151_req_1); -- 
    convTranspose_cp_element_group_384: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_384"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(382) & convTranspose_CP_39_elements(383);
      gj_convTranspose_cp_element_group_384 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(384), clk => clk, reset => reset); --
    end block;
    -- CP-element group 385:  merge  transition  place  bypass 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	381 
    -- CP-element group 385: 	384 
    -- CP-element group 385: successors 
    -- CP-element group 385: 	386 
    -- CP-element group 385:  members (2) 
      -- CP-element group 385: 	 branch_block_stmt_26/merge_stmt_1150_PhiAck/$entry
      -- CP-element group 385: 	 branch_block_stmt_26/merge_stmt_1150_PhiReqMerge
      -- 
    convTranspose_CP_39_elements(385) <= OrReduce(convTranspose_CP_39_elements(381) & convTranspose_CP_39_elements(384));
    -- CP-element group 386:  fork  transition  place  input  output  bypass 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	385 
    -- CP-element group 386: successors 
    -- CP-element group 386: 	312 
    -- CP-element group 386: 	313 
    -- CP-element group 386: 	315 
    -- CP-element group 386: 	317 
    -- CP-element group 386: 	319 
    -- CP-element group 386: 	321 
    -- CP-element group 386: 	323 
    -- CP-element group 386: 	325 
    -- CP-element group 386: 	327 
    -- CP-element group 386: 	329 
    -- CP-element group 386: 	331 
    -- CP-element group 386: 	333 
    -- CP-element group 386:  members (53) 
      -- CP-element group 386: 	 branch_block_stmt_26/merge_stmt_1150__exit__
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278__entry__
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/$entry
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/addr_of_1164_update_start_
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/array_obj_ref_1163_index_resized_1
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/array_obj_ref_1163_index_scaled_1
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/array_obj_ref_1163_index_computed_1
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/array_obj_ref_1163_index_resize_1/$entry
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/array_obj_ref_1163_index_resize_1/$exit
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/array_obj_ref_1163_index_resize_1/index_resize_req
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/array_obj_ref_1163_index_resize_1/index_resize_ack
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/array_obj_ref_1163_index_scale_1/$entry
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/array_obj_ref_1163_index_scale_1/$exit
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/array_obj_ref_1163_index_scale_1/scale_rename_req
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/array_obj_ref_1163_index_scale_1/scale_rename_ack
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/array_obj_ref_1163_final_index_sum_regn_update_start
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/array_obj_ref_1163_final_index_sum_regn_Sample/$entry
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/array_obj_ref_1163_final_index_sum_regn_Sample/req
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/array_obj_ref_1163_final_index_sum_regn_Update/$entry
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/array_obj_ref_1163_final_index_sum_regn_Update/req
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/addr_of_1164_complete/$entry
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/addr_of_1164_complete/req
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/ptr_deref_1168_update_start_
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/ptr_deref_1168_Update/$entry
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/ptr_deref_1168_Update/word_access_complete/$entry
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/ptr_deref_1168_Update/word_access_complete/word_0/$entry
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/ptr_deref_1168_Update/word_access_complete/word_0/cr
      -- CP-element group 386: 	 branch_block_stmt_26/merge_stmt_1150_PhiAck/phi_stmt_1151_ack
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1172_update_start_
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1172_Update/$entry
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1172_Update/cr
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1182_update_start_
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1182_Update/$entry
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1182_Update/cr
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1192_update_start_
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1192_Update/$entry
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1192_Update/cr
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1202_update_start_
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1202_Update/$entry
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1202_Update/cr
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1212_update_start_
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1212_Update/$entry
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1212_Update/cr
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1222_update_start_
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1222_Update/$entry
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1222_Update/cr
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1232_update_start_
      -- CP-element group 386: 	 branch_block_stmt_26/merge_stmt_1150_PhiAck/$exit
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1232_Update/$entry
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1232_Update/cr
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1242_update_start_
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1242_Update/$entry
      -- CP-element group 386: 	 branch_block_stmt_26/assign_stmt_1165_to_assign_stmt_1278/type_cast_1242_Update/cr
      -- 
    phi_stmt_1151_ack_3022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 386_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1151_ack_0, ack => convTranspose_CP_39_elements(386)); -- 
    req_2423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(386), ack => array_obj_ref_1163_index_offset_req_0); -- 
    req_2428_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2428_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(386), ack => array_obj_ref_1163_index_offset_req_1); -- 
    req_2443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(386), ack => addr_of_1164_final_reg_req_1); -- 
    cr_2488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(386), ack => ptr_deref_1168_load_0_req_1); -- 
    cr_2507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(386), ack => type_cast_1172_inst_req_1); -- 
    cr_2521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(386), ack => type_cast_1182_inst_req_1); -- 
    cr_2535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(386), ack => type_cast_1192_inst_req_1); -- 
    cr_2549_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2549_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(386), ack => type_cast_1202_inst_req_1); -- 
    cr_2563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(386), ack => type_cast_1212_inst_req_1); -- 
    cr_2577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(386), ack => type_cast_1222_inst_req_1); -- 
    cr_2591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(386), ack => type_cast_1232_inst_req_1); -- 
    cr_2605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(386), ack => type_cast_1242_inst_req_1); -- 
    -- CP-element group 387:  merge  transition  place  bypass 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	309 
    -- CP-element group 387: 	358 
    -- CP-element group 387: successors 
    -- CP-element group 387:  members (16) 
      -- CP-element group 387: 	 branch_block_stmt_26/branch_block_stmt_26__exit__
      -- CP-element group 387: 	 $exit
      -- CP-element group 387: 	 branch_block_stmt_26/$exit
      -- CP-element group 387: 	 branch_block_stmt_26/merge_stmt_1287__exit__
      -- CP-element group 387: 	 branch_block_stmt_26/return__
      -- CP-element group 387: 	 branch_block_stmt_26/merge_stmt_1289__exit__
      -- CP-element group 387: 	 branch_block_stmt_26/merge_stmt_1289_PhiAck/$exit
      -- CP-element group 387: 	 branch_block_stmt_26/merge_stmt_1289_PhiAck/dummy
      -- CP-element group 387: 	 branch_block_stmt_26/merge_stmt_1289_PhiAck/$entry
      -- CP-element group 387: 	 branch_block_stmt_26/merge_stmt_1289_PhiReqMerge
      -- CP-element group 387: 	 branch_block_stmt_26/return___PhiReq/$exit
      -- CP-element group 387: 	 branch_block_stmt_26/return___PhiReq/$entry
      -- CP-element group 387: 	 branch_block_stmt_26/merge_stmt_1287_PhiAck/dummy
      -- CP-element group 387: 	 branch_block_stmt_26/merge_stmt_1287_PhiAck/$exit
      -- CP-element group 387: 	 branch_block_stmt_26/merge_stmt_1287_PhiAck/$entry
      -- CP-element group 387: 	 branch_block_stmt_26/merge_stmt_1287_PhiReqMerge
      -- 
    convTranspose_CP_39_elements(387) <= OrReduce(convTranspose_CP_39_elements(309) & convTranspose_CP_39_elements(358));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar468_908_resized : std_logic_vector(13 downto 0);
    signal R_indvar468_908_scaled : std_logic_vector(13 downto 0);
    signal R_indvar482_664_resized : std_logic_vector(10 downto 0);
    signal R_indvar482_664_scaled : std_logic_vector(10 downto 0);
    signal R_indvar498_457_resized : std_logic_vector(13 downto 0);
    signal R_indvar498_457_scaled : std_logic_vector(13 downto 0);
    signal R_indvar_1162_resized : std_logic_vector(13 downto 0);
    signal R_indvar_1162_scaled : std_logic_vector(13 downto 0);
    signal add108_304 : std_logic_vector(15 downto 0);
    signal add117_329 : std_logic_vector(15 downto 0);
    signal add126_354 : std_logic_vector(15 downto 0);
    signal add12_76 : std_logic_vector(15 downto 0);
    signal add135_379 : std_logic_vector(15 downto 0);
    signal add150_485 : std_logic_vector(63 downto 0);
    signal add156_503 : std_logic_vector(63 downto 0);
    signal add162_521 : std_logic_vector(63 downto 0);
    signal add168_539 : std_logic_vector(63 downto 0);
    signal add174_557 : std_logic_vector(63 downto 0);
    signal add180_575 : std_logic_vector(63 downto 0);
    signal add186_593 : std_logic_vector(63 downto 0);
    signal add206_692 : std_logic_vector(63 downto 0);
    signal add212_710 : std_logic_vector(63 downto 0);
    signal add218_728 : std_logic_vector(63 downto 0);
    signal add21_101 : std_logic_vector(15 downto 0);
    signal add224_746 : std_logic_vector(63 downto 0);
    signal add230_764 : std_logic_vector(63 downto 0);
    signal add236_782 : std_logic_vector(63 downto 0);
    signal add242_800 : std_logic_vector(63 downto 0);
    signal add30_126 : std_logic_vector(15 downto 0);
    signal add39_151 : std_logic_vector(15 downto 0);
    signal add48_176 : std_logic_vector(15 downto 0);
    signal add57_201 : std_logic_vector(15 downto 0);
    signal add99_279 : std_logic_vector(15 downto 0);
    signal add_51 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1163_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1163_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1163_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1163_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1163_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1163_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_458_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_458_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_458_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_458_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_458_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_458_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_665_constant_part_of_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_665_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_665_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_665_offset_scale_factor_1 : std_logic_vector(10 downto 0);
    signal array_obj_ref_665_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_665_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_909_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_909_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_909_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_909_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_909_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_909_root_address : std_logic_vector(13 downto 0);
    signal arrayidx246_667 : std_logic_vector(31 downto 0);
    signal arrayidx269_911 : std_logic_vector(31 downto 0);
    signal arrayidx375_1165 : std_logic_vector(31 downto 0);
    signal arrayidx_460 : std_logic_vector(31 downto 0);
    signal call101_282 : std_logic_vector(7 downto 0);
    signal call106_295 : std_logic_vector(7 downto 0);
    signal call10_67 : std_logic_vector(7 downto 0);
    signal call110_307 : std_logic_vector(7 downto 0);
    signal call115_320 : std_logic_vector(7 downto 0);
    signal call119_332 : std_logic_vector(7 downto 0);
    signal call124_345 : std_logic_vector(7 downto 0);
    signal call128_357 : std_logic_vector(7 downto 0);
    signal call133_370 : std_logic_vector(7 downto 0);
    signal call143_463 : std_logic_vector(7 downto 0);
    signal call147_476 : std_logic_vector(7 downto 0);
    signal call14_79 : std_logic_vector(7 downto 0);
    signal call153_494 : std_logic_vector(7 downto 0);
    signal call159_512 : std_logic_vector(7 downto 0);
    signal call165_530 : std_logic_vector(7 downto 0);
    signal call171_548 : std_logic_vector(7 downto 0);
    signal call177_566 : std_logic_vector(7 downto 0);
    signal call183_584 : std_logic_vector(7 downto 0);
    signal call199_670 : std_logic_vector(7 downto 0);
    signal call19_92 : std_logic_vector(7 downto 0);
    signal call203_683 : std_logic_vector(7 downto 0);
    signal call209_701 : std_logic_vector(7 downto 0);
    signal call215_719 : std_logic_vector(7 downto 0);
    signal call221_737 : std_logic_vector(7 downto 0);
    signal call227_755 : std_logic_vector(7 downto 0);
    signal call233_773 : std_logic_vector(7 downto 0);
    signal call239_791 : std_logic_vector(7 downto 0);
    signal call23_104 : std_logic_vector(7 downto 0);
    signal call275_939 : std_logic_vector(63 downto 0);
    signal call28_117 : std_logic_vector(7 downto 0);
    signal call295_994 : std_logic_vector(15 downto 0);
    signal call297_997 : std_logic_vector(63 downto 0);
    signal call2_42 : std_logic_vector(7 downto 0);
    signal call32_129 : std_logic_vector(7 downto 0);
    signal call37_142 : std_logic_vector(7 downto 0);
    signal call41_154 : std_logic_vector(7 downto 0);
    signal call46_167 : std_logic_vector(7 downto 0);
    signal call50_179 : std_logic_vector(7 downto 0);
    signal call55_192 : std_logic_vector(7 downto 0);
    signal call5_54 : std_logic_vector(7 downto 0);
    signal call92_257 : std_logic_vector(7 downto 0);
    signal call97_270 : std_logic_vector(7 downto 0);
    signal call_29 : std_logic_vector(7 downto 0);
    signal cmp194452_401 : std_logic_vector(0 downto 0);
    signal cmp264448_852 : std_logic_vector(0 downto 0);
    signal cmp456_386 : std_logic_vector(0 downto 0);
    signal conv104_286 : std_logic_vector(15 downto 0);
    signal conv107_299 : std_logic_vector(15 downto 0);
    signal conv113_311 : std_logic_vector(15 downto 0);
    signal conv116_324 : std_logic_vector(15 downto 0);
    signal conv11_71 : std_logic_vector(15 downto 0);
    signal conv122_336 : std_logic_vector(15 downto 0);
    signal conv125_349 : std_logic_vector(15 downto 0);
    signal conv131_361 : std_logic_vector(15 downto 0);
    signal conv134_374 : std_logic_vector(15 downto 0);
    signal conv144_467 : std_logic_vector(63 downto 0);
    signal conv149_480 : std_logic_vector(63 downto 0);
    signal conv155_498 : std_logic_vector(63 downto 0);
    signal conv161_516 : std_logic_vector(63 downto 0);
    signal conv167_534 : std_logic_vector(63 downto 0);
    signal conv173_552 : std_logic_vector(63 downto 0);
    signal conv179_570 : std_logic_vector(63 downto 0);
    signal conv17_83 : std_logic_vector(15 downto 0);
    signal conv185_588 : std_logic_vector(63 downto 0);
    signal conv1_33 : std_logic_vector(15 downto 0);
    signal conv200_674 : std_logic_vector(63 downto 0);
    signal conv205_687 : std_logic_vector(63 downto 0);
    signal conv20_96 : std_logic_vector(15 downto 0);
    signal conv211_705 : std_logic_vector(63 downto 0);
    signal conv217_723 : std_logic_vector(63 downto 0);
    signal conv223_741 : std_logic_vector(63 downto 0);
    signal conv229_759 : std_logic_vector(63 downto 0);
    signal conv235_777 : std_logic_vector(63 downto 0);
    signal conv241_795 : std_logic_vector(63 downto 0);
    signal conv253_828 : std_logic_vector(31 downto 0);
    signal conv255_832 : std_logic_vector(31 downto 0);
    signal conv258_836 : std_logic_vector(31 downto 0);
    signal conv26_108 : std_logic_vector(15 downto 0);
    signal conv276_945 : std_logic_vector(63 downto 0);
    signal conv298_1002 : std_logic_vector(63 downto 0);
    signal conv29_121 : std_logic_vector(15 downto 0);
    signal conv304_1011 : std_logic_vector(7 downto 0);
    signal conv310_1021 : std_logic_vector(7 downto 0);
    signal conv316_1031 : std_logic_vector(7 downto 0);
    signal conv322_1041 : std_logic_vector(7 downto 0);
    signal conv328_1051 : std_logic_vector(7 downto 0);
    signal conv334_1061 : std_logic_vector(7 downto 0);
    signal conv340_1071 : std_logic_vector(7 downto 0);
    signal conv346_1081 : std_logic_vector(7 downto 0);
    signal conv35_133 : std_logic_vector(15 downto 0);
    signal conv380_1173 : std_logic_vector(7 downto 0);
    signal conv386_1183 : std_logic_vector(7 downto 0);
    signal conv38_146 : std_logic_vector(15 downto 0);
    signal conv392_1193 : std_logic_vector(7 downto 0);
    signal conv398_1203 : std_logic_vector(7 downto 0);
    signal conv3_46 : std_logic_vector(15 downto 0);
    signal conv404_1213 : std_logic_vector(7 downto 0);
    signal conv410_1223 : std_logic_vector(7 downto 0);
    signal conv416_1233 : std_logic_vector(7 downto 0);
    signal conv422_1243 : std_logic_vector(7 downto 0);
    signal conv44_158 : std_logic_vector(15 downto 0);
    signal conv47_171 : std_logic_vector(15 downto 0);
    signal conv53_183 : std_logic_vector(15 downto 0);
    signal conv56_196 : std_logic_vector(15 downto 0);
    signal conv61_205 : std_logic_vector(31 downto 0);
    signal conv63_209 : std_logic_vector(31 downto 0);
    signal conv65_213 : std_logic_vector(31 downto 0);
    signal conv82_227 : std_logic_vector(31 downto 0);
    signal conv84_231 : std_logic_vector(31 downto 0);
    signal conv87_235 : std_logic_vector(31 downto 0);
    signal conv8_58 : std_logic_vector(15 downto 0);
    signal conv90_239 : std_logic_vector(31 downto 0);
    signal conv95_261 : std_logic_vector(15 downto 0);
    signal conv98_274 : std_logic_vector(15 downto 0);
    signal exitcond1_1278 : std_logic_vector(0 downto 0);
    signal exitcond2_815 : std_logic_vector(0 downto 0);
    signal exitcond3_608 : std_logic_vector(0 downto 0);
    signal exitcond_927 : std_logic_vector(0 downto 0);
    signal iNsTr_108_1135 : std_logic_vector(63 downto 0);
    signal iNsTr_25_430 : std_logic_vector(63 downto 0);
    signal iNsTr_38_637 : std_logic_vector(63 downto 0);
    signal iNsTr_52_881 : std_logic_vector(63 downto 0);
    signal indvar468_897 : std_logic_vector(63 downto 0);
    signal indvar482_653 : std_logic_vector(63 downto 0);
    signal indvar498_446 : std_logic_vector(63 downto 0);
    signal indvar_1151 : std_logic_vector(63 downto 0);
    signal indvarx_xnext469_922 : std_logic_vector(63 downto 0);
    signal indvarx_xnext483_810 : std_logic_vector(63 downto 0);
    signal indvarx_xnext499_603 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1273 : std_logic_vector(63 downto 0);
    signal mul256_841 : std_logic_vector(31 downto 0);
    signal mul259_846 : std_logic_vector(31 downto 0);
    signal mul66_223 : std_logic_vector(31 downto 0);
    signal mul85_244 : std_logic_vector(31 downto 0);
    signal mul88_249 : std_logic_vector(31 downto 0);
    signal mul91_254 : std_logic_vector(31 downto 0);
    signal mul_218 : std_logic_vector(31 downto 0);
    signal ptr_deref_1168_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1168_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1168_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1168_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1168_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_595_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_595_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_595_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_595_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_595_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_595_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_802_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_802_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_802_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_802_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_802_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_802_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_913_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_913_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_913_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_913_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_913_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_913_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl105_292 : std_logic_vector(15 downto 0);
    signal shl114_317 : std_logic_vector(15 downto 0);
    signal shl123_342 : std_logic_vector(15 downto 0);
    signal shl132_367 : std_logic_vector(15 downto 0);
    signal shl146_473 : std_logic_vector(63 downto 0);
    signal shl152_491 : std_logic_vector(63 downto 0);
    signal shl158_509 : std_logic_vector(63 downto 0);
    signal shl164_527 : std_logic_vector(63 downto 0);
    signal shl170_545 : std_logic_vector(63 downto 0);
    signal shl176_563 : std_logic_vector(63 downto 0);
    signal shl182_581 : std_logic_vector(63 downto 0);
    signal shl18_89 : std_logic_vector(15 downto 0);
    signal shl202_680 : std_logic_vector(63 downto 0);
    signal shl208_698 : std_logic_vector(63 downto 0);
    signal shl214_716 : std_logic_vector(63 downto 0);
    signal shl220_734 : std_logic_vector(63 downto 0);
    signal shl226_752 : std_logic_vector(63 downto 0);
    signal shl232_770 : std_logic_vector(63 downto 0);
    signal shl238_788 : std_logic_vector(63 downto 0);
    signal shl27_114 : std_logic_vector(15 downto 0);
    signal shl36_139 : std_logic_vector(15 downto 0);
    signal shl45_164 : std_logic_vector(15 downto 0);
    signal shl54_189 : std_logic_vector(15 downto 0);
    signal shl96_267 : std_logic_vector(15 downto 0);
    signal shl9_64 : std_logic_vector(15 downto 0);
    signal shl_39 : std_logic_vector(15 downto 0);
    signal shr307_1017 : std_logic_vector(63 downto 0);
    signal shr313_1027 : std_logic_vector(63 downto 0);
    signal shr319_1037 : std_logic_vector(63 downto 0);
    signal shr325_1047 : std_logic_vector(63 downto 0);
    signal shr331_1057 : std_logic_vector(63 downto 0);
    signal shr337_1067 : std_logic_vector(63 downto 0);
    signal shr343_1077 : std_logic_vector(63 downto 0);
    signal shr383_1179 : std_logic_vector(63 downto 0);
    signal shr389_1189 : std_logic_vector(63 downto 0);
    signal shr395_1199 : std_logic_vector(63 downto 0);
    signal shr401_1209 : std_logic_vector(63 downto 0);
    signal shr407_1219 : std_logic_vector(63 downto 0);
    signal shr413_1229 : std_logic_vector(63 downto 0);
    signal shr419_1239 : std_logic_vector(63 downto 0);
    signal sub_1007 : std_logic_vector(63 downto 0);
    signal tmp376_1169 : std_logic_vector(63 downto 0);
    signal tmp463_1119 : std_logic_vector(31 downto 0);
    signal tmp463x_xop_1131 : std_logic_vector(31 downto 0);
    signal tmp464_1125 : std_logic_vector(0 downto 0);
    signal tmp467_1148 : std_logic_vector(63 downto 0);
    signal tmp475_865 : std_logic_vector(31 downto 0);
    signal tmp475x_xop_877 : std_logic_vector(31 downto 0);
    signal tmp476_871 : std_logic_vector(0 downto 0);
    signal tmp480_894 : std_logic_vector(63 downto 0);
    signal tmp491_621 : std_logic_vector(31 downto 0);
    signal tmp491x_xop_633 : std_logic_vector(31 downto 0);
    signal tmp492_627 : std_logic_vector(0 downto 0);
    signal tmp496_650 : std_logic_vector(63 downto 0);
    signal tmp505_414 : std_logic_vector(31 downto 0);
    signal tmp505x_xop_426 : std_logic_vector(31 downto 0);
    signal tmp506_420 : std_logic_vector(0 downto 0);
    signal tmp510_443 : std_logic_vector(63 downto 0);
    signal type_cast_1000_wire : std_logic_vector(63 downto 0);
    signal type_cast_1015_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1025_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1035_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1045_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1055_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1065_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1075_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1117_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1123_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1129_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_112_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1139_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1146_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1155_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1157_wire : std_logic_vector(63 downto 0);
    signal type_cast_1177_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1187_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1197_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1207_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1217_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1227_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1237_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1271_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_137_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_162_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_187_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_265_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_290_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_315_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_340_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_365_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_37_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_383_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_399_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_412_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_418_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_424_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_434_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_441_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_450_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_452_wire : std_logic_vector(63 downto 0);
    signal type_cast_471_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_489_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_507_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_525_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_543_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_561_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_579_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_601_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_619_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_625_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_62_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_631_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_641_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_648_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_657_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_659_wire : std_logic_vector(63 downto 0);
    signal type_cast_678_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_696_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_714_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_732_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_750_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_768_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_786_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_808_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_850_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_863_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_869_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_875_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_87_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_885_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_892_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_901_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_903_wire : std_logic_vector(63 downto 0);
    signal type_cast_915_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_920_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_943_wire : std_logic_vector(63 downto 0);
    signal type_cast_976_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_980_wire_constant : std_logic_vector(15 downto 0);
    signal xx_xop512_887 : std_logic_vector(63 downto 0);
    signal xx_xop513_643 : std_logic_vector(63 downto 0);
    signal xx_xop514_436 : std_logic_vector(63 downto 0);
    signal xx_xop_1141 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1163_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1163_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1163_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1163_resized_base_address <= "00000000000000";
    array_obj_ref_458_constant_part_of_offset <= "00000000000000";
    array_obj_ref_458_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_458_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_458_resized_base_address <= "00000000000000";
    array_obj_ref_665_constant_part_of_offset <= "00000100010";
    array_obj_ref_665_offset_scale_factor_0 <= "10000000000";
    array_obj_ref_665_offset_scale_factor_1 <= "00000000001";
    array_obj_ref_665_resized_base_address <= "00000000000";
    array_obj_ref_909_constant_part_of_offset <= "00000000000000";
    array_obj_ref_909_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_909_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_909_resized_base_address <= "00000000000000";
    ptr_deref_1168_word_offset_0 <= "00000000000000";
    ptr_deref_595_word_offset_0 <= "00000000000000";
    ptr_deref_802_word_offset_0 <= "00000000000";
    ptr_deref_913_word_offset_0 <= "00000000000000";
    type_cast_1015_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1025_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1035_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1045_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1055_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1065_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1075_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1117_wire_constant <= "00000000000000000000000000000010";
    type_cast_1123_wire_constant <= "00000000000000000000000000000001";
    type_cast_1129_wire_constant <= "11111111111111111111111111111111";
    type_cast_112_wire_constant <= "0000000000001000";
    type_cast_1139_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1146_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1155_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1177_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1187_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1197_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1207_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1217_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1227_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1237_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1271_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_137_wire_constant <= "0000000000001000";
    type_cast_162_wire_constant <= "0000000000001000";
    type_cast_187_wire_constant <= "0000000000001000";
    type_cast_265_wire_constant <= "0000000000001000";
    type_cast_290_wire_constant <= "0000000000001000";
    type_cast_315_wire_constant <= "0000000000001000";
    type_cast_340_wire_constant <= "0000000000001000";
    type_cast_365_wire_constant <= "0000000000001000";
    type_cast_37_wire_constant <= "0000000000001000";
    type_cast_383_wire_constant <= "00000000000000000000000000000011";
    type_cast_399_wire_constant <= "00000000000000000000000000000011";
    type_cast_412_wire_constant <= "00000000000000000000000000000010";
    type_cast_418_wire_constant <= "00000000000000000000000000000001";
    type_cast_424_wire_constant <= "11111111111111111111111111111111";
    type_cast_434_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_441_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_450_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_471_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_489_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_507_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_525_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_543_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_561_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_579_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_601_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_619_wire_constant <= "00000000000000000000000000000010";
    type_cast_625_wire_constant <= "00000000000000000000000000000001";
    type_cast_62_wire_constant <= "0000000000001000";
    type_cast_631_wire_constant <= "11111111111111111111111111111111";
    type_cast_641_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_648_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_657_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_678_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_696_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_714_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_732_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_750_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_768_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_786_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_808_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_850_wire_constant <= "00000000000000000000000000000011";
    type_cast_863_wire_constant <= "00000000000000000000000000000010";
    type_cast_869_wire_constant <= "00000000000000000000000000000001";
    type_cast_875_wire_constant <= "11111111111111111111111111111111";
    type_cast_87_wire_constant <= "0000000000001000";
    type_cast_885_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_892_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_901_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_915_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_920_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_976_wire_constant <= "0000000000000000";
    type_cast_980_wire_constant <= "0000000000000000";
    phi_stmt_1151: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1155_wire_constant & type_cast_1157_wire;
      req <= phi_stmt_1151_req_0 & phi_stmt_1151_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1151",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1151_ack_0,
          idata => idata,
          odata => indvar_1151,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1151
    phi_stmt_446: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_450_wire_constant & type_cast_452_wire;
      req <= phi_stmt_446_req_0 & phi_stmt_446_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_446",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_446_ack_0,
          idata => idata,
          odata => indvar498_446,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_446
    phi_stmt_653: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_657_wire_constant & type_cast_659_wire;
      req <= phi_stmt_653_req_0 & phi_stmt_653_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_653",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_653_ack_0,
          idata => idata,
          odata => indvar482_653,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_653
    phi_stmt_897: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_901_wire_constant & type_cast_903_wire;
      req <= phi_stmt_897_req_0 & phi_stmt_897_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_897",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_897_ack_0,
          idata => idata,
          odata => indvar468_897,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_897
    -- flow-through select operator MUX_1147_inst
    tmp467_1148 <= xx_xop_1141 when (tmp464_1125(0) /=  '0') else type_cast_1146_wire_constant;
    -- flow-through select operator MUX_442_inst
    tmp510_443 <= xx_xop514_436 when (tmp506_420(0) /=  '0') else type_cast_441_wire_constant;
    -- flow-through select operator MUX_649_inst
    tmp496_650 <= xx_xop513_643 when (tmp492_627(0) /=  '0') else type_cast_648_wire_constant;
    -- flow-through select operator MUX_893_inst
    tmp480_894 <= xx_xop512_887 when (tmp476_871(0) /=  '0') else type_cast_892_wire_constant;
    addr_of_1164_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1164_final_reg_req_0;
      addr_of_1164_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1164_final_reg_req_1;
      addr_of_1164_final_reg_ack_1<= rack(0);
      addr_of_1164_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1164_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1163_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx375_1165,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_459_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_459_final_reg_req_0;
      addr_of_459_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_459_final_reg_req_1;
      addr_of_459_final_reg_ack_1<= rack(0);
      addr_of_459_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_459_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_458_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_460,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_666_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_666_final_reg_req_0;
      addr_of_666_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_666_final_reg_req_1;
      addr_of_666_final_reg_ack_1<= rack(0);
      addr_of_666_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_666_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 11,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_665_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx246_667,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_910_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_910_final_reg_req_0;
      addr_of_910_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_910_final_reg_req_1;
      addr_of_910_final_reg_ack_1<= rack(0);
      addr_of_910_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_910_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_909_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx269_911,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1001_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1001_inst_req_0;
      type_cast_1001_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1001_inst_req_1;
      type_cast_1001_inst_ack_1<= rack(0);
      type_cast_1001_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1001_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1000_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv298_1002,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1010_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1010_inst_req_0;
      type_cast_1010_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1010_inst_req_1;
      type_cast_1010_inst_ack_1<= rack(0);
      type_cast_1010_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1010_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub_1007,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv304_1011,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1020_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1020_inst_req_0;
      type_cast_1020_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1020_inst_req_1;
      type_cast_1020_inst_ack_1<= rack(0);
      type_cast_1020_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1020_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr307_1017,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv310_1021,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1030_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1030_inst_req_0;
      type_cast_1030_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1030_inst_req_1;
      type_cast_1030_inst_ack_1<= rack(0);
      type_cast_1030_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1030_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr313_1027,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv316_1031,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1040_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1040_inst_req_0;
      type_cast_1040_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1040_inst_req_1;
      type_cast_1040_inst_ack_1<= rack(0);
      type_cast_1040_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1040_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr319_1037,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv322_1041,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1050_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1050_inst_req_0;
      type_cast_1050_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1050_inst_req_1;
      type_cast_1050_inst_ack_1<= rack(0);
      type_cast_1050_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1050_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr325_1047,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv328_1051,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1060_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1060_inst_req_0;
      type_cast_1060_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1060_inst_req_1;
      type_cast_1060_inst_ack_1<= rack(0);
      type_cast_1060_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1060_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr331_1057,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv334_1061,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1070_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1070_inst_req_0;
      type_cast_1070_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1070_inst_req_1;
      type_cast_1070_inst_ack_1<= rack(0);
      type_cast_1070_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1070_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr337_1067,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv340_1071,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_107_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_107_inst_req_0;
      type_cast_107_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_107_inst_req_1;
      type_cast_107_inst_ack_1<= rack(0);
      type_cast_107_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_107_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call23_104,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv26_108,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1080_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1080_inst_req_0;
      type_cast_1080_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1080_inst_req_1;
      type_cast_1080_inst_ack_1<= rack(0);
      type_cast_1080_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1080_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr343_1077,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv346_1081,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1134_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1134_inst_req_0;
      type_cast_1134_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1134_inst_req_1;
      type_cast_1134_inst_ack_1<= rack(0);
      type_cast_1134_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1134_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp463x_xop_1131,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_108_1135,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1157_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1157_inst_req_0;
      type_cast_1157_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1157_inst_req_1;
      type_cast_1157_inst_ack_1<= rack(0);
      type_cast_1157_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1157_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1273,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1157_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1172_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1172_inst_req_0;
      type_cast_1172_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1172_inst_req_1;
      type_cast_1172_inst_ack_1<= rack(0);
      type_cast_1172_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1172_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp376_1169,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv380_1173,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1182_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1182_inst_req_0;
      type_cast_1182_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1182_inst_req_1;
      type_cast_1182_inst_ack_1<= rack(0);
      type_cast_1182_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1182_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr383_1179,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv386_1183,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1192_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1192_inst_req_0;
      type_cast_1192_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1192_inst_req_1;
      type_cast_1192_inst_ack_1<= rack(0);
      type_cast_1192_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1192_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr389_1189,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv392_1193,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1202_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1202_inst_req_0;
      type_cast_1202_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1202_inst_req_1;
      type_cast_1202_inst_ack_1<= rack(0);
      type_cast_1202_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1202_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr395_1199,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv398_1203,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_120_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_120_inst_req_0;
      type_cast_120_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_120_inst_req_1;
      type_cast_120_inst_ack_1<= rack(0);
      type_cast_120_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_120_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call28_117,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_121,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1212_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1212_inst_req_0;
      type_cast_1212_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1212_inst_req_1;
      type_cast_1212_inst_ack_1<= rack(0);
      type_cast_1212_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1212_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr401_1209,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv404_1213,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1222_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1222_inst_req_0;
      type_cast_1222_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1222_inst_req_1;
      type_cast_1222_inst_ack_1<= rack(0);
      type_cast_1222_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1222_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr407_1219,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv410_1223,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1232_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1232_inst_req_0;
      type_cast_1232_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1232_inst_req_1;
      type_cast_1232_inst_ack_1<= rack(0);
      type_cast_1232_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1232_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr413_1229,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv416_1233,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1242_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1242_inst_req_0;
      type_cast_1242_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1242_inst_req_1;
      type_cast_1242_inst_ack_1<= rack(0);
      type_cast_1242_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1242_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr419_1239,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv422_1243,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_132_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_132_inst_req_0;
      type_cast_132_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_132_inst_req_1;
      type_cast_132_inst_ack_1<= rack(0);
      type_cast_132_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_132_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call32_129,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv35_133,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_145_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_145_inst_req_0;
      type_cast_145_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_145_inst_req_1;
      type_cast_145_inst_ack_1<= rack(0);
      type_cast_145_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_145_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call37_142,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_146,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_157_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_157_inst_req_0;
      type_cast_157_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_157_inst_req_1;
      type_cast_157_inst_ack_1<= rack(0);
      type_cast_157_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_157_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_154,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_158,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_170_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_170_inst_req_0;
      type_cast_170_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_170_inst_req_1;
      type_cast_170_inst_ack_1<= rack(0);
      type_cast_170_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_170_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_167,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv47_171,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_182_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_182_inst_req_0;
      type_cast_182_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_182_inst_req_1;
      type_cast_182_inst_ack_1<= rack(0);
      type_cast_182_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_182_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call50_179,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv53_183,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_195_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_195_inst_req_0;
      type_cast_195_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_195_inst_req_1;
      type_cast_195_inst_ack_1<= rack(0);
      type_cast_195_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_195_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call55_192,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_196,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_204_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_204_inst_req_0;
      type_cast_204_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_204_inst_req_1;
      type_cast_204_inst_ack_1<= rack(0);
      type_cast_204_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_204_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_51,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv61_205,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_208_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_208_inst_req_0;
      type_cast_208_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_208_inst_req_1;
      type_cast_208_inst_ack_1<= rack(0);
      type_cast_208_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_208_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add12_76,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv63_209,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_212_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_212_inst_req_0;
      type_cast_212_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_212_inst_req_1;
      type_cast_212_inst_ack_1<= rack(0);
      type_cast_212_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_212_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add21_101,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_213,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_226_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_226_inst_req_0;
      type_cast_226_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_226_inst_req_1;
      type_cast_226_inst_ack_1<= rack(0);
      type_cast_226_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_226_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add30_126,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv82_227,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_230_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_230_inst_req_0;
      type_cast_230_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_230_inst_req_1;
      type_cast_230_inst_ack_1<= rack(0);
      type_cast_230_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_230_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add39_151,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv84_231,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_234_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_234_inst_req_0;
      type_cast_234_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_234_inst_req_1;
      type_cast_234_inst_ack_1<= rack(0);
      type_cast_234_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_234_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add48_176,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv87_235,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_238_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_238_inst_req_0;
      type_cast_238_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_238_inst_req_1;
      type_cast_238_inst_ack_1<= rack(0);
      type_cast_238_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_238_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add57_201,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_239,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_260_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_260_inst_req_0;
      type_cast_260_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_260_inst_req_1;
      type_cast_260_inst_ack_1<= rack(0);
      type_cast_260_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_260_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call92_257,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_261,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_273_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_273_inst_req_0;
      type_cast_273_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_273_inst_req_1;
      type_cast_273_inst_ack_1<= rack(0);
      type_cast_273_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_273_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call97_270,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv98_274,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_285_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_285_inst_req_0;
      type_cast_285_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_285_inst_req_1;
      type_cast_285_inst_ack_1<= rack(0);
      type_cast_285_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_285_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call101_282,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv104_286,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_298_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_298_inst_req_0;
      type_cast_298_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_298_inst_req_1;
      type_cast_298_inst_ack_1<= rack(0);
      type_cast_298_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_298_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call106_295,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv107_299,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_310_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_310_inst_req_0;
      type_cast_310_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_310_inst_req_1;
      type_cast_310_inst_ack_1<= rack(0);
      type_cast_310_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_310_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call110_307,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv113_311,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_323_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_323_inst_req_0;
      type_cast_323_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_323_inst_req_1;
      type_cast_323_inst_ack_1<= rack(0);
      type_cast_323_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_323_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call115_320,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv116_324,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_32_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_32_inst_req_0;
      type_cast_32_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_32_inst_req_1;
      type_cast_32_inst_ack_1<= rack(0);
      type_cast_32_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_32_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_29,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1_33,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_335_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_335_inst_req_0;
      type_cast_335_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_335_inst_req_1;
      type_cast_335_inst_ack_1<= rack(0);
      type_cast_335_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_335_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call119_332,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv122_336,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_348_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_348_inst_req_0;
      type_cast_348_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_348_inst_req_1;
      type_cast_348_inst_ack_1<= rack(0);
      type_cast_348_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_348_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call124_345,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv125_349,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_360_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_360_inst_req_0;
      type_cast_360_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_360_inst_req_1;
      type_cast_360_inst_ack_1<= rack(0);
      type_cast_360_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_360_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call128_357,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv131_361,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_373_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_373_inst_req_0;
      type_cast_373_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_373_inst_req_1;
      type_cast_373_inst_ack_1<= rack(0);
      type_cast_373_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_373_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call133_370,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv134_374,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_429_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_429_inst_req_0;
      type_cast_429_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_429_inst_req_1;
      type_cast_429_inst_ack_1<= rack(0);
      type_cast_429_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_429_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp505x_xop_426,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_25_430,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_452_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_452_inst_req_0;
      type_cast_452_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_452_inst_req_1;
      type_cast_452_inst_ack_1<= rack(0);
      type_cast_452_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_452_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext499_603,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_452_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_45_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_45_inst_req_0;
      type_cast_45_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_45_inst_req_1;
      type_cast_45_inst_ack_1<= rack(0);
      type_cast_45_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_45_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_42,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_46,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_466_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_466_inst_req_0;
      type_cast_466_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_466_inst_req_1;
      type_cast_466_inst_ack_1<= rack(0);
      type_cast_466_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_466_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call143_463,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv144_467,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_479_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_479_inst_req_0;
      type_cast_479_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_479_inst_req_1;
      type_cast_479_inst_ack_1<= rack(0);
      type_cast_479_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_479_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call147_476,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv149_480,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_497_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_497_inst_req_0;
      type_cast_497_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_497_inst_req_1;
      type_cast_497_inst_ack_1<= rack(0);
      type_cast_497_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_497_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call153_494,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv155_498,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_515_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_515_inst_req_0;
      type_cast_515_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_515_inst_req_1;
      type_cast_515_inst_ack_1<= rack(0);
      type_cast_515_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_515_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call159_512,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv161_516,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_533_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_533_inst_req_0;
      type_cast_533_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_533_inst_req_1;
      type_cast_533_inst_ack_1<= rack(0);
      type_cast_533_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_533_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call165_530,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv167_534,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_551_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_551_inst_req_0;
      type_cast_551_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_551_inst_req_1;
      type_cast_551_inst_ack_1<= rack(0);
      type_cast_551_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_551_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call171_548,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv173_552,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_569_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_569_inst_req_0;
      type_cast_569_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_569_inst_req_1;
      type_cast_569_inst_ack_1<= rack(0);
      type_cast_569_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_569_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call177_566,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv179_570,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_57_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_57_inst_req_0;
      type_cast_57_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_57_inst_req_1;
      type_cast_57_inst_ack_1<= rack(0);
      type_cast_57_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_57_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_54,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv8_58,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_587_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_587_inst_req_0;
      type_cast_587_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_587_inst_req_1;
      type_cast_587_inst_ack_1<= rack(0);
      type_cast_587_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_587_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call183_584,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv185_588,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_636_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_636_inst_req_0;
      type_cast_636_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_636_inst_req_1;
      type_cast_636_inst_ack_1<= rack(0);
      type_cast_636_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_636_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp491x_xop_633,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_38_637,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_659_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_659_inst_req_0;
      type_cast_659_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_659_inst_req_1;
      type_cast_659_inst_ack_1<= rack(0);
      type_cast_659_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_659_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext483_810,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_659_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_673_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_673_inst_req_0;
      type_cast_673_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_673_inst_req_1;
      type_cast_673_inst_ack_1<= rack(0);
      type_cast_673_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_673_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call199_670,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv200_674,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_686_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_686_inst_req_0;
      type_cast_686_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_686_inst_req_1;
      type_cast_686_inst_ack_1<= rack(0);
      type_cast_686_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_686_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call203_683,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv205_687,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_704_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_704_inst_req_0;
      type_cast_704_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_704_inst_req_1;
      type_cast_704_inst_ack_1<= rack(0);
      type_cast_704_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_704_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call209_701,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv211_705,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_70_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_70_inst_req_0;
      type_cast_70_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_70_inst_req_1;
      type_cast_70_inst_ack_1<= rack(0);
      type_cast_70_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_70_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call10_67,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv11_71,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_722_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_722_inst_req_0;
      type_cast_722_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_722_inst_req_1;
      type_cast_722_inst_ack_1<= rack(0);
      type_cast_722_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_722_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call215_719,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv217_723,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_740_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_740_inst_req_0;
      type_cast_740_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_740_inst_req_1;
      type_cast_740_inst_ack_1<= rack(0);
      type_cast_740_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_740_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call221_737,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv223_741,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_758_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_758_inst_req_0;
      type_cast_758_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_758_inst_req_1;
      type_cast_758_inst_ack_1<= rack(0);
      type_cast_758_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_758_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call227_755,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv229_759,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_776_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_776_inst_req_0;
      type_cast_776_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_776_inst_req_1;
      type_cast_776_inst_ack_1<= rack(0);
      type_cast_776_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_776_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call233_773,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv235_777,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_794_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_794_inst_req_0;
      type_cast_794_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_794_inst_req_1;
      type_cast_794_inst_ack_1<= rack(0);
      type_cast_794_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_794_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call239_791,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv241_795,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_827_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_827_inst_req_0;
      type_cast_827_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_827_inst_req_1;
      type_cast_827_inst_ack_1<= rack(0);
      type_cast_827_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_827_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add117_329,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv253_828,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_82_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_82_inst_req_0;
      type_cast_82_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_82_inst_req_1;
      type_cast_82_inst_ack_1<= rack(0);
      type_cast_82_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_82_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call14_79,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_83,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_831_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_831_inst_req_0;
      type_cast_831_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_831_inst_req_1;
      type_cast_831_inst_ack_1<= rack(0);
      type_cast_831_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_831_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add126_354,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv255_832,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_835_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_835_inst_req_0;
      type_cast_835_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_835_inst_req_1;
      type_cast_835_inst_ack_1<= rack(0);
      type_cast_835_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_835_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add135_379,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv258_836,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_880_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_880_inst_req_0;
      type_cast_880_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_880_inst_req_1;
      type_cast_880_inst_ack_1<= rack(0);
      type_cast_880_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_880_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp475x_xop_877,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_52_881,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_903_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_903_inst_req_0;
      type_cast_903_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_903_inst_req_1;
      type_cast_903_inst_ack_1<= rack(0);
      type_cast_903_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_903_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext469_922,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_903_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_944_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_944_inst_req_0;
      type_cast_944_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_944_inst_req_1;
      type_cast_944_inst_ack_1<= rack(0);
      type_cast_944_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_944_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_943_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv276_945,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_95_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_95_inst_req_0;
      type_cast_95_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_95_inst_req_1;
      type_cast_95_inst_ack_1<= rack(0);
      type_cast_95_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_95_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call19_92,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv20_96,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1163_index_1_rename
    process(R_indvar_1162_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_1162_resized;
      ov(13 downto 0) := iv;
      R_indvar_1162_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1163_index_1_resize
    process(indvar_1151) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_1151;
      ov := iv(13 downto 0);
      R_indvar_1162_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1163_root_address_inst
    process(array_obj_ref_1163_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1163_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1163_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_458_index_1_rename
    process(R_indvar498_457_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar498_457_resized;
      ov(13 downto 0) := iv;
      R_indvar498_457_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_458_index_1_resize
    process(indvar498_446) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar498_446;
      ov := iv(13 downto 0);
      R_indvar498_457_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_458_root_address_inst
    process(array_obj_ref_458_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_458_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_458_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_665_index_1_rename
    process(R_indvar482_664_resized) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar482_664_resized;
      ov(10 downto 0) := iv;
      R_indvar482_664_scaled <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_665_index_1_resize
    process(indvar482_653) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar482_653;
      ov := iv(10 downto 0);
      R_indvar482_664_resized <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_665_root_address_inst
    process(array_obj_ref_665_final_offset) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_665_final_offset;
      ov(10 downto 0) := iv;
      array_obj_ref_665_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_909_index_1_rename
    process(R_indvar468_908_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar468_908_resized;
      ov(13 downto 0) := iv;
      R_indvar468_908_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_909_index_1_resize
    process(indvar468_897) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar468_897;
      ov := iv(13 downto 0);
      R_indvar468_908_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_909_root_address_inst
    process(array_obj_ref_909_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_909_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_909_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1168_addr_0
    process(ptr_deref_1168_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1168_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1168_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1168_base_resize
    process(arrayidx375_1165) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx375_1165;
      ov := iv(13 downto 0);
      ptr_deref_1168_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1168_gather_scatter
    process(ptr_deref_1168_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1168_data_0;
      ov(63 downto 0) := iv;
      tmp376_1169 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1168_root_address_inst
    process(ptr_deref_1168_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1168_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1168_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_595_addr_0
    process(ptr_deref_595_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_595_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_595_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_595_base_resize
    process(arrayidx_460) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_460;
      ov := iv(13 downto 0);
      ptr_deref_595_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_595_gather_scatter
    process(add186_593) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add186_593;
      ov(63 downto 0) := iv;
      ptr_deref_595_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_595_root_address_inst
    process(ptr_deref_595_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_595_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_595_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_802_addr_0
    process(ptr_deref_802_root_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_802_root_address;
      ov(10 downto 0) := iv;
      ptr_deref_802_word_address_0 <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_802_base_resize
    process(arrayidx246_667) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx246_667;
      ov := iv(10 downto 0);
      ptr_deref_802_resized_base_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_802_gather_scatter
    process(add242_800) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add242_800;
      ov(63 downto 0) := iv;
      ptr_deref_802_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_802_root_address_inst
    process(ptr_deref_802_resized_base_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_802_resized_base_address;
      ov(10 downto 0) := iv;
      ptr_deref_802_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_913_addr_0
    process(ptr_deref_913_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_913_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_913_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_913_base_resize
    process(arrayidx269_911) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx269_911;
      ov := iv(13 downto 0);
      ptr_deref_913_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_913_gather_scatter
    process(type_cast_915_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_915_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_913_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_913_root_address_inst
    process(ptr_deref_913_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_913_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_913_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1107_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp264448_852;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1107_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1107_branch_req_0,
          ack0 => if_stmt_1107_branch_ack_0,
          ack1 => if_stmt_1107_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1279_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_1278;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1279_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1279_branch_req_0,
          ack0 => if_stmt_1279_branch_ack_0,
          ack1 => if_stmt_1279_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_387_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp456_386;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_387_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_387_branch_req_0,
          ack0 => if_stmt_387_branch_ack_0,
          ack1 => if_stmt_387_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_402_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp194452_401;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_402_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_402_branch_req_0,
          ack0 => if_stmt_402_branch_ack_0,
          ack1 => if_stmt_402_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_609_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond3_608;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_609_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_609_branch_req_0,
          ack0 => if_stmt_609_branch_ack_0,
          ack1 => if_stmt_609_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_816_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond2_815;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_816_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_816_branch_req_0,
          ack0 => if_stmt_816_branch_ack_0,
          ack1 => if_stmt_816_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_853_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp264448_852;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_853_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_853_branch_req_0,
          ack0 => if_stmt_853_branch_ack_0,
          ack1 => if_stmt_853_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_928_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_927;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_928_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_928_branch_req_0,
          ack0 => if_stmt_928_branch_ack_0,
          ack1 => if_stmt_928_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_1130_inst
    process(tmp463_1119) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp463_1119, type_cast_1129_wire_constant, tmp_var);
      tmp463x_xop_1131 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_425_inst
    process(tmp505_414) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp505_414, type_cast_424_wire_constant, tmp_var);
      tmp505x_xop_426 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_632_inst
    process(tmp491_621) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp491_621, type_cast_631_wire_constant, tmp_var);
      tmp491x_xop_633 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_876_inst
    process(tmp475_865) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp475_865, type_cast_875_wire_constant, tmp_var);
      tmp475x_xop_877 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1140_inst
    process(iNsTr_108_1135) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_108_1135, type_cast_1139_wire_constant, tmp_var);
      xx_xop_1141 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1272_inst
    process(indvar_1151) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1151, type_cast_1271_wire_constant, tmp_var);
      indvarx_xnext_1273 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_435_inst
    process(iNsTr_25_430) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_25_430, type_cast_434_wire_constant, tmp_var);
      xx_xop514_436 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_602_inst
    process(indvar498_446) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar498_446, type_cast_601_wire_constant, tmp_var);
      indvarx_xnext499_603 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_642_inst
    process(iNsTr_38_637) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_38_637, type_cast_641_wire_constant, tmp_var);
      xx_xop513_643 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_809_inst
    process(indvar482_653) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar482_653, type_cast_808_wire_constant, tmp_var);
      indvarx_xnext483_810 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_886_inst
    process(iNsTr_52_881) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_52_881, type_cast_885_wire_constant, tmp_var);
      xx_xop512_887 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_921_inst
    process(indvar468_897) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar468_897, type_cast_920_wire_constant, tmp_var);
      indvarx_xnext469_922 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1277_inst
    process(indvarx_xnext_1273, tmp467_1148) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1273, tmp467_1148, tmp_var);
      exitcond1_1278 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_607_inst
    process(indvarx_xnext499_603, tmp510_443) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext499_603, tmp510_443, tmp_var);
      exitcond3_608 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_814_inst
    process(indvarx_xnext483_810, tmp496_650) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext483_810, tmp496_650, tmp_var);
      exitcond2_815 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_926_inst
    process(indvarx_xnext469_922, tmp480_894) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext469_922, tmp480_894, tmp_var);
      exitcond_927 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1118_inst
    process(mul259_846) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul259_846, type_cast_1117_wire_constant, tmp_var);
      tmp463_1119 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_413_inst
    process(mul66_223) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_223, type_cast_412_wire_constant, tmp_var);
      tmp505_414 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_620_inst
    process(mul91_254) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul91_254, type_cast_619_wire_constant, tmp_var);
      tmp491_621 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_864_inst
    process(mul259_846) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul259_846, type_cast_863_wire_constant, tmp_var);
      tmp475_865 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1016_inst
    process(sub_1007) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1007, type_cast_1015_wire_constant, tmp_var);
      shr307_1017 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1026_inst
    process(sub_1007) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1007, type_cast_1025_wire_constant, tmp_var);
      shr313_1027 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1036_inst
    process(sub_1007) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1007, type_cast_1035_wire_constant, tmp_var);
      shr319_1037 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1046_inst
    process(sub_1007) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1007, type_cast_1045_wire_constant, tmp_var);
      shr325_1047 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1056_inst
    process(sub_1007) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1007, type_cast_1055_wire_constant, tmp_var);
      shr331_1057 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1066_inst
    process(sub_1007) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1007, type_cast_1065_wire_constant, tmp_var);
      shr337_1067 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1076_inst
    process(sub_1007) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1007, type_cast_1075_wire_constant, tmp_var);
      shr343_1077 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1178_inst
    process(tmp376_1169) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp376_1169, type_cast_1177_wire_constant, tmp_var);
      shr383_1179 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1188_inst
    process(tmp376_1169) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp376_1169, type_cast_1187_wire_constant, tmp_var);
      shr389_1189 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1198_inst
    process(tmp376_1169) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp376_1169, type_cast_1197_wire_constant, tmp_var);
      shr395_1199 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1208_inst
    process(tmp376_1169) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp376_1169, type_cast_1207_wire_constant, tmp_var);
      shr401_1209 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1218_inst
    process(tmp376_1169) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp376_1169, type_cast_1217_wire_constant, tmp_var);
      shr407_1219 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1228_inst
    process(tmp376_1169) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp376_1169, type_cast_1227_wire_constant, tmp_var);
      shr413_1229 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1238_inst
    process(tmp376_1169) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp376_1169, type_cast_1237_wire_constant, tmp_var);
      shr419_1239 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_217_inst
    process(conv63_209, conv61_205) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv63_209, conv61_205, tmp_var);
      mul_218 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_222_inst
    process(mul_218, conv65_213) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_218, conv65_213, tmp_var);
      mul66_223 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_243_inst
    process(conv84_231, conv82_227) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv84_231, conv82_227, tmp_var);
      mul85_244 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_248_inst
    process(mul85_244, conv87_235) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul85_244, conv87_235, tmp_var);
      mul88_249 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_253_inst
    process(mul88_249, conv90_239) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul88_249, conv90_239, tmp_var);
      mul91_254 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_840_inst
    process(conv255_832, conv253_828) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv255_832, conv253_828, tmp_var);
      mul256_841 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_845_inst
    process(mul256_841, conv258_836) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul256_841, conv258_836, tmp_var);
      mul259_846 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_100_inst
    process(shl18_89, conv20_96) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl18_89, conv20_96, tmp_var);
      add21_101 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_125_inst
    process(shl27_114, conv29_121) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl27_114, conv29_121, tmp_var);
      add30_126 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_150_inst
    process(shl36_139, conv38_146) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl36_139, conv38_146, tmp_var);
      add39_151 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_175_inst
    process(shl45_164, conv47_171) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl45_164, conv47_171, tmp_var);
      add48_176 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_200_inst
    process(shl54_189, conv56_196) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl54_189, conv56_196, tmp_var);
      add57_201 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_278_inst
    process(shl96_267, conv98_274) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl96_267, conv98_274, tmp_var);
      add99_279 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_303_inst
    process(shl105_292, conv107_299) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl105_292, conv107_299, tmp_var);
      add108_304 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_328_inst
    process(shl114_317, conv116_324) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl114_317, conv116_324, tmp_var);
      add117_329 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_353_inst
    process(shl123_342, conv125_349) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl123_342, conv125_349, tmp_var);
      add126_354 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_378_inst
    process(shl132_367, conv134_374) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl132_367, conv134_374, tmp_var);
      add135_379 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_50_inst
    process(shl_39, conv3_46) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_39, conv3_46, tmp_var);
      add_51 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_75_inst
    process(shl9_64, conv11_71) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl9_64, conv11_71, tmp_var);
      add12_76 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_484_inst
    process(shl146_473, conv149_480) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl146_473, conv149_480, tmp_var);
      add150_485 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_502_inst
    process(shl152_491, conv155_498) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl152_491, conv155_498, tmp_var);
      add156_503 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_520_inst
    process(shl158_509, conv161_516) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl158_509, conv161_516, tmp_var);
      add162_521 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_538_inst
    process(shl164_527, conv167_534) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl164_527, conv167_534, tmp_var);
      add168_539 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_556_inst
    process(shl170_545, conv173_552) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl170_545, conv173_552, tmp_var);
      add174_557 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_574_inst
    process(shl176_563, conv179_570) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl176_563, conv179_570, tmp_var);
      add180_575 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_592_inst
    process(shl182_581, conv185_588) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl182_581, conv185_588, tmp_var);
      add186_593 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_691_inst
    process(shl202_680, conv205_687) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl202_680, conv205_687, tmp_var);
      add206_692 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_709_inst
    process(shl208_698, conv211_705) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl208_698, conv211_705, tmp_var);
      add212_710 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_727_inst
    process(shl214_716, conv217_723) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl214_716, conv217_723, tmp_var);
      add218_728 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_745_inst
    process(shl220_734, conv223_741) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl220_734, conv223_741, tmp_var);
      add224_746 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_763_inst
    process(shl226_752, conv229_759) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl226_752, conv229_759, tmp_var);
      add230_764 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_781_inst
    process(shl232_770, conv235_777) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl232_770, conv235_777, tmp_var);
      add236_782 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_799_inst
    process(shl238_788, conv241_795) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl238_788, conv241_795, tmp_var);
      add242_800 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_113_inst
    process(conv26_108) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv26_108, type_cast_112_wire_constant, tmp_var);
      shl27_114 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_138_inst
    process(conv35_133) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv35_133, type_cast_137_wire_constant, tmp_var);
      shl36_139 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_163_inst
    process(conv44_158) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv44_158, type_cast_162_wire_constant, tmp_var);
      shl45_164 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_188_inst
    process(conv53_183) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv53_183, type_cast_187_wire_constant, tmp_var);
      shl54_189 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_266_inst
    process(conv95_261) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv95_261, type_cast_265_wire_constant, tmp_var);
      shl96_267 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_291_inst
    process(conv104_286) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv104_286, type_cast_290_wire_constant, tmp_var);
      shl105_292 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_316_inst
    process(conv113_311) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv113_311, type_cast_315_wire_constant, tmp_var);
      shl114_317 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_341_inst
    process(conv122_336) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv122_336, type_cast_340_wire_constant, tmp_var);
      shl123_342 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_366_inst
    process(conv131_361) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv131_361, type_cast_365_wire_constant, tmp_var);
      shl132_367 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_38_inst
    process(conv1_33) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1_33, type_cast_37_wire_constant, tmp_var);
      shl_39 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_63_inst
    process(conv8_58) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv8_58, type_cast_62_wire_constant, tmp_var);
      shl9_64 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_88_inst
    process(conv17_83) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv17_83, type_cast_87_wire_constant, tmp_var);
      shl18_89 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_472_inst
    process(conv144_467) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv144_467, type_cast_471_wire_constant, tmp_var);
      shl146_473 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_490_inst
    process(add150_485) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add150_485, type_cast_489_wire_constant, tmp_var);
      shl152_491 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_508_inst
    process(add156_503) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add156_503, type_cast_507_wire_constant, tmp_var);
      shl158_509 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_526_inst
    process(add162_521) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add162_521, type_cast_525_wire_constant, tmp_var);
      shl164_527 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_544_inst
    process(add168_539) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add168_539, type_cast_543_wire_constant, tmp_var);
      shl170_545 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_562_inst
    process(add174_557) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add174_557, type_cast_561_wire_constant, tmp_var);
      shl176_563 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_580_inst
    process(add180_575) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add180_575, type_cast_579_wire_constant, tmp_var);
      shl182_581 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_679_inst
    process(conv200_674) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv200_674, type_cast_678_wire_constant, tmp_var);
      shl202_680 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_697_inst
    process(add206_692) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add206_692, type_cast_696_wire_constant, tmp_var);
      shl208_698 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_715_inst
    process(add212_710) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add212_710, type_cast_714_wire_constant, tmp_var);
      shl214_716 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_733_inst
    process(add218_728) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add218_728, type_cast_732_wire_constant, tmp_var);
      shl220_734 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_751_inst
    process(add224_746) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add224_746, type_cast_750_wire_constant, tmp_var);
      shl226_752 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_769_inst
    process(add230_764) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add230_764, type_cast_768_wire_constant, tmp_var);
      shl232_770 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_787_inst
    process(add236_782) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add236_782, type_cast_786_wire_constant, tmp_var);
      shl238_788 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_1006_inst
    process(conv298_1002, conv276_945) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv298_1002, conv276_945, tmp_var);
      sub_1007 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1124_inst
    process(tmp463_1119) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp463_1119, type_cast_1123_wire_constant, tmp_var);
      tmp464_1125 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_384_inst
    process(mul66_223) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul66_223, type_cast_383_wire_constant, tmp_var);
      cmp456_386 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_400_inst
    process(mul91_254) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul91_254, type_cast_399_wire_constant, tmp_var);
      cmp194452_401 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_419_inst
    process(tmp505_414) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp505_414, type_cast_418_wire_constant, tmp_var);
      tmp506_420 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_626_inst
    process(tmp491_621) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp491_621, type_cast_625_wire_constant, tmp_var);
      tmp492_627 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_851_inst
    process(mul259_846) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul259_846, type_cast_850_wire_constant, tmp_var);
      cmp264448_852 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_870_inst
    process(tmp475_865) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp475_865, type_cast_869_wire_constant, tmp_var);
      tmp476_871 <= tmp_var; --
    end process;
    -- shared split operator group (101) : array_obj_ref_1163_index_offset 
    ApIntAdd_group_101: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_1162_scaled;
      array_obj_ref_1163_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1163_index_offset_req_0;
      array_obj_ref_1163_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1163_index_offset_req_1;
      array_obj_ref_1163_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_101_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_101_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_101",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 101
    -- shared split operator group (102) : array_obj_ref_458_index_offset 
    ApIntAdd_group_102: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar498_457_scaled;
      array_obj_ref_458_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_458_index_offset_req_0;
      array_obj_ref_458_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_458_index_offset_req_1;
      array_obj_ref_458_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_102_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_102_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_102",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 102
    -- shared split operator group (103) : array_obj_ref_665_index_offset 
    ApIntAdd_group_103: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar482_664_scaled;
      array_obj_ref_665_final_offset <= data_out(10 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_665_index_offset_req_0;
      array_obj_ref_665_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_665_index_offset_req_1;
      array_obj_ref_665_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_103_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_103_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_103",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000100010",
          constant_width => 11,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 103
    -- shared split operator group (104) : array_obj_ref_909_index_offset 
    ApIntAdd_group_104: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar468_908_scaled;
      array_obj_ref_909_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_909_index_offset_req_0;
      array_obj_ref_909_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_909_index_offset_req_1;
      array_obj_ref_909_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_104_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_104_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_104",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 104
    -- unary operator type_cast_1000_inst
    process(call297_997) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call297_997, tmp_var);
      type_cast_1000_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_943_inst
    process(call275_939) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call275_939, tmp_var);
      type_cast_943_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_1168_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1168_load_0_req_0;
      ptr_deref_1168_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1168_load_0_req_1;
      ptr_deref_1168_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1168_word_address_0;
      ptr_deref_1168_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(13 downto 0),
          mtag => memory_space_3_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(63 downto 0),
          mtag => memory_space_3_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_595_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_595_store_0_req_0;
      ptr_deref_595_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_595_store_0_req_1;
      ptr_deref_595_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_595_word_address_0;
      data_in <= ptr_deref_595_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_802_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(10 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_802_store_0_req_0;
      ptr_deref_802_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_802_store_0_req_1;
      ptr_deref_802_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_802_word_address_0;
      data_in <= ptr_deref_802_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 11,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(10 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_913_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_913_store_0_req_0;
      ptr_deref_913_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_913_store_0_req_1;
      ptr_deref_913_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_913_word_address_0;
      data_in <= ptr_deref_913_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared inport operator group (0) : RPIPE_Block0_done_993_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block0_done_993_inst_req_0;
      RPIPE_Block0_done_993_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block0_done_993_inst_req_1;
      RPIPE_Block0_done_993_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call295_994 <= data_out(15 downto 0);
      Block0_done_read_0_gI: SplitGuardInterface generic map(name => "Block0_done_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_done_read_0: InputPortRevised -- 
        generic map ( name => "Block0_done_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_done_pipe_read_req(0),
          oack => Block0_done_pipe_read_ack(0),
          odata => Block0_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_ConvTranspose_input_pipe_565_inst RPIPE_ConvTranspose_input_pipe_547_inst RPIPE_ConvTranspose_input_pipe_583_inst RPIPE_ConvTranspose_input_pipe_475_inst RPIPE_ConvTranspose_input_pipe_529_inst RPIPE_ConvTranspose_input_pipe_669_inst RPIPE_ConvTranspose_input_pipe_462_inst RPIPE_ConvTranspose_input_pipe_682_inst RPIPE_ConvTranspose_input_pipe_700_inst RPIPE_ConvTranspose_input_pipe_511_inst RPIPE_ConvTranspose_input_pipe_718_inst RPIPE_ConvTranspose_input_pipe_736_inst RPIPE_ConvTranspose_input_pipe_754_inst RPIPE_ConvTranspose_input_pipe_493_inst RPIPE_ConvTranspose_input_pipe_772_inst RPIPE_ConvTranspose_input_pipe_790_inst RPIPE_ConvTranspose_input_pipe_28_inst RPIPE_ConvTranspose_input_pipe_41_inst RPIPE_ConvTranspose_input_pipe_53_inst RPIPE_ConvTranspose_input_pipe_66_inst RPIPE_ConvTranspose_input_pipe_78_inst RPIPE_ConvTranspose_input_pipe_91_inst RPIPE_ConvTranspose_input_pipe_103_inst RPIPE_ConvTranspose_input_pipe_116_inst RPIPE_ConvTranspose_input_pipe_128_inst RPIPE_ConvTranspose_input_pipe_141_inst RPIPE_ConvTranspose_input_pipe_153_inst RPIPE_ConvTranspose_input_pipe_166_inst RPIPE_ConvTranspose_input_pipe_178_inst RPIPE_ConvTranspose_input_pipe_191_inst RPIPE_ConvTranspose_input_pipe_256_inst RPIPE_ConvTranspose_input_pipe_269_inst RPIPE_ConvTranspose_input_pipe_281_inst RPIPE_ConvTranspose_input_pipe_294_inst RPIPE_ConvTranspose_input_pipe_306_inst RPIPE_ConvTranspose_input_pipe_319_inst RPIPE_ConvTranspose_input_pipe_331_inst RPIPE_ConvTranspose_input_pipe_344_inst RPIPE_ConvTranspose_input_pipe_356_inst RPIPE_ConvTranspose_input_pipe_369_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(319 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 39 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 39 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 39 downto 0);
      signal guard_vector : std_logic_vector( 39 downto 0);
      constant outBUFs : IntegerArray(39 downto 0) := (39 => 1, 38 => 1, 37 => 1, 36 => 1, 35 => 1, 34 => 1, 33 => 1, 32 => 1, 31 => 1, 30 => 1, 29 => 1, 28 => 1, 27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(39 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false, 28 => false, 29 => false, 30 => false, 31 => false, 32 => false, 33 => false, 34 => false, 35 => false, 36 => false, 37 => false, 38 => false, 39 => false);
      constant guardBuffering: IntegerArray(39 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2, 28 => 2, 29 => 2, 30 => 2, 31 => 2, 32 => 2, 33 => 2, 34 => 2, 35 => 2, 36 => 2, 37 => 2, 38 => 2, 39 => 2);
      -- 
    begin -- 
      reqL_unguarded(39) <= RPIPE_ConvTranspose_input_pipe_565_inst_req_0;
      reqL_unguarded(38) <= RPIPE_ConvTranspose_input_pipe_547_inst_req_0;
      reqL_unguarded(37) <= RPIPE_ConvTranspose_input_pipe_583_inst_req_0;
      reqL_unguarded(36) <= RPIPE_ConvTranspose_input_pipe_475_inst_req_0;
      reqL_unguarded(35) <= RPIPE_ConvTranspose_input_pipe_529_inst_req_0;
      reqL_unguarded(34) <= RPIPE_ConvTranspose_input_pipe_669_inst_req_0;
      reqL_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_462_inst_req_0;
      reqL_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_682_inst_req_0;
      reqL_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_700_inst_req_0;
      reqL_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_511_inst_req_0;
      reqL_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_718_inst_req_0;
      reqL_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_736_inst_req_0;
      reqL_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_754_inst_req_0;
      reqL_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_493_inst_req_0;
      reqL_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_772_inst_req_0;
      reqL_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_790_inst_req_0;
      reqL_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_28_inst_req_0;
      reqL_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_41_inst_req_0;
      reqL_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_53_inst_req_0;
      reqL_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_66_inst_req_0;
      reqL_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_78_inst_req_0;
      reqL_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_91_inst_req_0;
      reqL_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_103_inst_req_0;
      reqL_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_116_inst_req_0;
      reqL_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_128_inst_req_0;
      reqL_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_141_inst_req_0;
      reqL_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_153_inst_req_0;
      reqL_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_166_inst_req_0;
      reqL_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_178_inst_req_0;
      reqL_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_191_inst_req_0;
      reqL_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_256_inst_req_0;
      reqL_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_269_inst_req_0;
      reqL_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_281_inst_req_0;
      reqL_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_294_inst_req_0;
      reqL_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_306_inst_req_0;
      reqL_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_319_inst_req_0;
      reqL_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_331_inst_req_0;
      reqL_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_344_inst_req_0;
      reqL_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_356_inst_req_0;
      reqL_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_369_inst_req_0;
      RPIPE_ConvTranspose_input_pipe_565_inst_ack_0 <= ackL_unguarded(39);
      RPIPE_ConvTranspose_input_pipe_547_inst_ack_0 <= ackL_unguarded(38);
      RPIPE_ConvTranspose_input_pipe_583_inst_ack_0 <= ackL_unguarded(37);
      RPIPE_ConvTranspose_input_pipe_475_inst_ack_0 <= ackL_unguarded(36);
      RPIPE_ConvTranspose_input_pipe_529_inst_ack_0 <= ackL_unguarded(35);
      RPIPE_ConvTranspose_input_pipe_669_inst_ack_0 <= ackL_unguarded(34);
      RPIPE_ConvTranspose_input_pipe_462_inst_ack_0 <= ackL_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_682_inst_ack_0 <= ackL_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_700_inst_ack_0 <= ackL_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_511_inst_ack_0 <= ackL_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_718_inst_ack_0 <= ackL_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_736_inst_ack_0 <= ackL_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_754_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_493_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_772_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_790_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_28_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_41_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_53_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_66_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_78_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_91_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_103_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_116_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_128_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_141_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_153_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_166_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_178_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_191_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_256_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_269_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_281_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_294_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_306_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_319_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_331_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_344_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_356_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_369_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(39) <= RPIPE_ConvTranspose_input_pipe_565_inst_req_1;
      reqR_unguarded(38) <= RPIPE_ConvTranspose_input_pipe_547_inst_req_1;
      reqR_unguarded(37) <= RPIPE_ConvTranspose_input_pipe_583_inst_req_1;
      reqR_unguarded(36) <= RPIPE_ConvTranspose_input_pipe_475_inst_req_1;
      reqR_unguarded(35) <= RPIPE_ConvTranspose_input_pipe_529_inst_req_1;
      reqR_unguarded(34) <= RPIPE_ConvTranspose_input_pipe_669_inst_req_1;
      reqR_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_462_inst_req_1;
      reqR_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_682_inst_req_1;
      reqR_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_700_inst_req_1;
      reqR_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_511_inst_req_1;
      reqR_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_718_inst_req_1;
      reqR_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_736_inst_req_1;
      reqR_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_754_inst_req_1;
      reqR_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_493_inst_req_1;
      reqR_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_772_inst_req_1;
      reqR_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_790_inst_req_1;
      reqR_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_28_inst_req_1;
      reqR_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_41_inst_req_1;
      reqR_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_53_inst_req_1;
      reqR_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_66_inst_req_1;
      reqR_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_78_inst_req_1;
      reqR_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_91_inst_req_1;
      reqR_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_103_inst_req_1;
      reqR_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_116_inst_req_1;
      reqR_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_128_inst_req_1;
      reqR_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_141_inst_req_1;
      reqR_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_153_inst_req_1;
      reqR_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_166_inst_req_1;
      reqR_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_178_inst_req_1;
      reqR_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_191_inst_req_1;
      reqR_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_256_inst_req_1;
      reqR_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_269_inst_req_1;
      reqR_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_281_inst_req_1;
      reqR_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_294_inst_req_1;
      reqR_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_306_inst_req_1;
      reqR_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_319_inst_req_1;
      reqR_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_331_inst_req_1;
      reqR_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_344_inst_req_1;
      reqR_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_356_inst_req_1;
      reqR_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_369_inst_req_1;
      RPIPE_ConvTranspose_input_pipe_565_inst_ack_1 <= ackR_unguarded(39);
      RPIPE_ConvTranspose_input_pipe_547_inst_ack_1 <= ackR_unguarded(38);
      RPIPE_ConvTranspose_input_pipe_583_inst_ack_1 <= ackR_unguarded(37);
      RPIPE_ConvTranspose_input_pipe_475_inst_ack_1 <= ackR_unguarded(36);
      RPIPE_ConvTranspose_input_pipe_529_inst_ack_1 <= ackR_unguarded(35);
      RPIPE_ConvTranspose_input_pipe_669_inst_ack_1 <= ackR_unguarded(34);
      RPIPE_ConvTranspose_input_pipe_462_inst_ack_1 <= ackR_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_682_inst_ack_1 <= ackR_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_700_inst_ack_1 <= ackR_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_511_inst_ack_1 <= ackR_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_718_inst_ack_1 <= ackR_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_736_inst_ack_1 <= ackR_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_754_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_493_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_772_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_790_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_28_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_41_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_53_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_66_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_78_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_91_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_103_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_116_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_128_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_141_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_153_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_166_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_178_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_191_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_256_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_269_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_281_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_294_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_306_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_319_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_331_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_344_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_356_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_369_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      guard_vector(34)  <=  '1';
      guard_vector(35)  <=  '1';
      guard_vector(36)  <=  '1';
      guard_vector(37)  <=  '1';
      guard_vector(38)  <=  '1';
      guard_vector(39)  <=  '1';
      call177_566 <= data_out(319 downto 312);
      call171_548 <= data_out(311 downto 304);
      call183_584 <= data_out(303 downto 296);
      call147_476 <= data_out(295 downto 288);
      call165_530 <= data_out(287 downto 280);
      call199_670 <= data_out(279 downto 272);
      call143_463 <= data_out(271 downto 264);
      call203_683 <= data_out(263 downto 256);
      call209_701 <= data_out(255 downto 248);
      call159_512 <= data_out(247 downto 240);
      call215_719 <= data_out(239 downto 232);
      call221_737 <= data_out(231 downto 224);
      call227_755 <= data_out(223 downto 216);
      call153_494 <= data_out(215 downto 208);
      call233_773 <= data_out(207 downto 200);
      call239_791 <= data_out(199 downto 192);
      call_29 <= data_out(191 downto 184);
      call2_42 <= data_out(183 downto 176);
      call5_54 <= data_out(175 downto 168);
      call10_67 <= data_out(167 downto 160);
      call14_79 <= data_out(159 downto 152);
      call19_92 <= data_out(151 downto 144);
      call23_104 <= data_out(143 downto 136);
      call28_117 <= data_out(135 downto 128);
      call32_129 <= data_out(127 downto 120);
      call37_142 <= data_out(119 downto 112);
      call41_154 <= data_out(111 downto 104);
      call46_167 <= data_out(103 downto 96);
      call50_179 <= data_out(95 downto 88);
      call55_192 <= data_out(87 downto 80);
      call92_257 <= data_out(79 downto 72);
      call97_270 <= data_out(71 downto 64);
      call101_282 <= data_out(63 downto 56);
      call106_295 <= data_out(55 downto 48);
      call110_307 <= data_out(47 downto 40);
      call115_320 <= data_out(39 downto 32);
      call119_332 <= data_out(31 downto 24);
      call124_345 <= data_out(23 downto 16);
      call128_357 <= data_out(15 downto 8);
      call133_370 <= data_out(7 downto 0);
      ConvTranspose_input_pipe_read_1_gI: SplitGuardInterface generic map(name => "ConvTranspose_input_pipe_read_1_gI", nreqs => 40, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_input_pipe_read_1: InputPortRevised -- 
        generic map ( name => "ConvTranspose_input_pipe_read_1", data_width => 8,  num_reqs => 40,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => ConvTranspose_input_pipe_pipe_read_req(0),
          oack => ConvTranspose_input_pipe_pipe_read_ack(0),
          odata => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared outport operator group (0) : WPIPE_Block0_start_965_inst WPIPE_Block0_start_962_inst WPIPE_Block0_start_985_inst WPIPE_Block0_start_959_inst WPIPE_Block0_start_968_inst WPIPE_Block0_start_971_inst WPIPE_Block0_start_988_inst WPIPE_Block0_start_974_inst WPIPE_Block0_start_978_inst WPIPE_Block0_start_982_inst WPIPE_Block0_start_953_inst WPIPE_Block0_start_956_inst WPIPE_Block0_start_950_inst WPIPE_Block0_start_947_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block0_start_965_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block0_start_962_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block0_start_985_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block0_start_959_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block0_start_968_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block0_start_971_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block0_start_988_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block0_start_974_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block0_start_978_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block0_start_982_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block0_start_953_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block0_start_956_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block0_start_950_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block0_start_947_inst_req_0;
      WPIPE_Block0_start_965_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block0_start_962_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block0_start_985_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block0_start_959_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block0_start_968_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block0_start_971_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block0_start_988_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block0_start_974_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block0_start_978_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block0_start_982_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block0_start_953_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block0_start_956_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block0_start_950_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block0_start_947_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block0_start_965_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block0_start_962_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block0_start_985_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block0_start_959_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block0_start_968_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block0_start_971_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block0_start_988_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block0_start_974_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block0_start_978_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block0_start_982_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block0_start_953_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block0_start_956_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block0_start_950_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block0_start_947_inst_req_1;
      WPIPE_Block0_start_965_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block0_start_962_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block0_start_985_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block0_start_959_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block0_start_968_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block0_start_971_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block0_start_988_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block0_start_974_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block0_start_978_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block0_start_982_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block0_start_953_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block0_start_956_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block0_start_950_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block0_start_947_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= add57_201 & add48_176 & add126_354 & add39_151 & add99_279 & add108_304 & add135_379 & type_cast_976_wire_constant & type_cast_980_wire_constant & add117_329 & add21_101 & add30_126 & add12_76 & add_51;
      Block0_start_write_0_gI: SplitGuardInterface generic map(name => "Block0_start_write_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_start_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_start_pipe_write_req(0),
          oack => Block0_start_pipe_write_ack(0),
          odata => Block0_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_ConvTranspose_output_pipe_1088_inst WPIPE_ConvTranspose_output_pipe_1091_inst WPIPE_ConvTranspose_output_pipe_1085_inst WPIPE_ConvTranspose_output_pipe_1097_inst WPIPE_ConvTranspose_output_pipe_1094_inst WPIPE_ConvTranspose_output_pipe_1082_inst WPIPE_ConvTranspose_output_pipe_1100_inst WPIPE_ConvTranspose_output_pipe_1103_inst WPIPE_ConvTranspose_output_pipe_1244_inst WPIPE_ConvTranspose_output_pipe_1247_inst WPIPE_ConvTranspose_output_pipe_1250_inst WPIPE_ConvTranspose_output_pipe_1253_inst WPIPE_ConvTranspose_output_pipe_1256_inst WPIPE_ConvTranspose_output_pipe_1259_inst WPIPE_ConvTranspose_output_pipe_1262_inst WPIPE_ConvTranspose_output_pipe_1265_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal sample_req, sample_ack : BooleanArray( 15 downto 0);
      signal update_req, update_ack : BooleanArray( 15 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 15 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 15 downto 0);
      signal guard_vector : std_logic_vector( 15 downto 0);
      constant inBUFs : IntegerArray(15 downto 0) := (15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(15 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false);
      constant guardBuffering: IntegerArray(15 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2);
      -- 
    begin -- 
      sample_req_unguarded(15) <= WPIPE_ConvTranspose_output_pipe_1088_inst_req_0;
      sample_req_unguarded(14) <= WPIPE_ConvTranspose_output_pipe_1091_inst_req_0;
      sample_req_unguarded(13) <= WPIPE_ConvTranspose_output_pipe_1085_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_ConvTranspose_output_pipe_1097_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_ConvTranspose_output_pipe_1094_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_ConvTranspose_output_pipe_1082_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_ConvTranspose_output_pipe_1100_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_ConvTranspose_output_pipe_1103_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1244_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1247_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1250_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1253_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1256_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1259_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1262_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1265_inst_req_0;
      WPIPE_ConvTranspose_output_pipe_1088_inst_ack_0 <= sample_ack_unguarded(15);
      WPIPE_ConvTranspose_output_pipe_1091_inst_ack_0 <= sample_ack_unguarded(14);
      WPIPE_ConvTranspose_output_pipe_1085_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_ConvTranspose_output_pipe_1097_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_ConvTranspose_output_pipe_1094_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_ConvTranspose_output_pipe_1082_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_ConvTranspose_output_pipe_1100_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_ConvTranspose_output_pipe_1103_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_ConvTranspose_output_pipe_1244_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1247_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1250_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1253_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1256_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1259_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1262_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1265_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(15) <= WPIPE_ConvTranspose_output_pipe_1088_inst_req_1;
      update_req_unguarded(14) <= WPIPE_ConvTranspose_output_pipe_1091_inst_req_1;
      update_req_unguarded(13) <= WPIPE_ConvTranspose_output_pipe_1085_inst_req_1;
      update_req_unguarded(12) <= WPIPE_ConvTranspose_output_pipe_1097_inst_req_1;
      update_req_unguarded(11) <= WPIPE_ConvTranspose_output_pipe_1094_inst_req_1;
      update_req_unguarded(10) <= WPIPE_ConvTranspose_output_pipe_1082_inst_req_1;
      update_req_unguarded(9) <= WPIPE_ConvTranspose_output_pipe_1100_inst_req_1;
      update_req_unguarded(8) <= WPIPE_ConvTranspose_output_pipe_1103_inst_req_1;
      update_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1244_inst_req_1;
      update_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1247_inst_req_1;
      update_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1250_inst_req_1;
      update_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1253_inst_req_1;
      update_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1256_inst_req_1;
      update_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1259_inst_req_1;
      update_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1262_inst_req_1;
      update_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1265_inst_req_1;
      WPIPE_ConvTranspose_output_pipe_1088_inst_ack_1 <= update_ack_unguarded(15);
      WPIPE_ConvTranspose_output_pipe_1091_inst_ack_1 <= update_ack_unguarded(14);
      WPIPE_ConvTranspose_output_pipe_1085_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_ConvTranspose_output_pipe_1097_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_ConvTranspose_output_pipe_1094_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_ConvTranspose_output_pipe_1082_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_ConvTranspose_output_pipe_1100_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_ConvTranspose_output_pipe_1103_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_ConvTranspose_output_pipe_1244_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1247_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1250_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1253_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1256_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1259_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1262_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1265_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      data_in <= conv334_1061 & conv328_1051 & conv340_1071 & conv316_1031 & conv322_1041 & conv346_1081 & conv310_1021 & conv304_1011 & conv422_1243 & conv416_1233 & conv410_1223 & conv404_1213 & conv398_1203 & conv392_1193 & conv386_1183 & conv380_1173;
      ConvTranspose_output_pipe_write_1_gI: SplitGuardInterface generic map(name => "ConvTranspose_output_pipe_write_1_gI", nreqs => 16, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_output_pipe_write_1: OutputPortRevised -- 
        generic map ( name => "ConvTranspose_output_pipe", data_width => 8, num_reqs => 16, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => ConvTranspose_output_pipe_pipe_write_req(0),
          oack => ConvTranspose_output_pipe_pipe_write_ack(0),
          odata => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_939_call call_stmt_997_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_939_call_req_0;
      reqL_unguarded(0) <= call_stmt_997_call_req_0;
      call_stmt_939_call_ack_0 <= ackL_unguarded(1);
      call_stmt_997_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_939_call_req_1;
      reqR_unguarded(0) <= call_stmt_997_call_req_1;
      call_stmt_939_call_ack_1 <= ackR_unguarded(1);
      call_stmt_997_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call275_939 <= data_out(127 downto 64);
      call297_997 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end convTranspose_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeA is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeA;
architecture convTransposeA_arch of convTransposeA is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeA_CP_3054_start: Boolean;
  signal convTransposeA_CP_3054_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_1339_inst_req_0 : boolean;
  signal type_cast_1380_inst_req_0 : boolean;
  signal type_cast_1380_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1347_inst_req_1 : boolean;
  signal type_cast_1326_inst_ack_1 : boolean;
  signal type_cast_1384_inst_ack_1 : boolean;
  signal type_cast_1392_inst_req_1 : boolean;
  signal type_cast_1326_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1347_inst_ack_1 : boolean;
  signal type_cast_1388_inst_ack_1 : boolean;
  signal type_cast_1472_inst_ack_0 : boolean;
  signal type_cast_1392_inst_ack_1 : boolean;
  signal type_cast_1339_inst_ack_0 : boolean;
  signal type_cast_1472_inst_req_1 : boolean;
  signal type_cast_1502_inst_req_0 : boolean;
  signal type_cast_1380_inst_req_1 : boolean;
  signal type_cast_1502_inst_req_1 : boolean;
  signal type_cast_1468_inst_ack_1 : boolean;
  signal type_cast_1339_inst_req_1 : boolean;
  signal type_cast_1339_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1350_inst_req_0 : boolean;
  signal type_cast_1380_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1347_inst_req_0 : boolean;
  signal type_cast_1384_inst_req_0 : boolean;
  signal type_cast_1502_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1350_inst_ack_0 : boolean;
  signal type_cast_1464_inst_req_1 : boolean;
  signal type_cast_1472_inst_req_0 : boolean;
  signal type_cast_1464_inst_ack_1 : boolean;
  signal type_cast_1472_inst_ack_1 : boolean;
  signal type_cast_1384_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1353_inst_req_0 : boolean;
  signal type_cast_1502_inst_ack_1 : boolean;
  signal type_cast_1468_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1335_inst_req_0 : boolean;
  signal type_cast_1392_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1353_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1347_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1350_inst_req_1 : boolean;
  signal type_cast_1392_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1353_inst_req_1 : boolean;
  signal type_cast_1388_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1335_inst_ack_0 : boolean;
  signal type_cast_1468_inst_req_1 : boolean;
  signal type_cast_1388_inst_ack_0 : boolean;
  signal type_cast_1464_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1350_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1353_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1335_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1335_inst_ack_1 : boolean;
  signal type_cast_1464_inst_ack_0 : boolean;
  signal type_cast_1384_inst_req_1 : boolean;
  signal type_cast_1468_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1295_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1295_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1295_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1295_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1298_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1298_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1298_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1298_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1301_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1301_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1301_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1301_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1304_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1304_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1304_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1304_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1307_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1307_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1307_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1307_inst_ack_1 : boolean;
  signal type_cast_1388_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1310_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1310_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1310_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1310_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1313_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1313_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1313_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1313_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1316_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1316_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1316_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1316_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1319_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1319_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1319_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1319_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1322_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1322_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1322_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1322_inst_ack_1 : boolean;
  signal type_cast_1326_inst_req_0 : boolean;
  signal type_cast_1326_inst_ack_0 : boolean;
  signal array_obj_ref_1508_index_offset_req_0 : boolean;
  signal array_obj_ref_1508_index_offset_ack_0 : boolean;
  signal array_obj_ref_1508_index_offset_req_1 : boolean;
  signal array_obj_ref_1508_index_offset_ack_1 : boolean;
  signal addr_of_1509_final_reg_req_0 : boolean;
  signal addr_of_1509_final_reg_ack_0 : boolean;
  signal addr_of_1509_final_reg_req_1 : boolean;
  signal addr_of_1509_final_reg_ack_1 : boolean;
  signal ptr_deref_1513_load_0_req_0 : boolean;
  signal ptr_deref_1513_load_0_ack_0 : boolean;
  signal ptr_deref_1513_load_0_req_1 : boolean;
  signal ptr_deref_1513_load_0_ack_1 : boolean;
  signal array_obj_ref_1531_index_offset_req_0 : boolean;
  signal array_obj_ref_1531_index_offset_ack_0 : boolean;
  signal array_obj_ref_1531_index_offset_req_1 : boolean;
  signal array_obj_ref_1531_index_offset_ack_1 : boolean;
  signal addr_of_1532_final_reg_req_0 : boolean;
  signal addr_of_1532_final_reg_ack_0 : boolean;
  signal addr_of_1532_final_reg_req_1 : boolean;
  signal addr_of_1532_final_reg_ack_1 : boolean;
  signal ptr_deref_1535_store_0_req_0 : boolean;
  signal ptr_deref_1535_store_0_ack_0 : boolean;
  signal ptr_deref_1535_store_0_req_1 : boolean;
  signal ptr_deref_1535_store_0_ack_1 : boolean;
  signal type_cast_1540_inst_req_0 : boolean;
  signal type_cast_1540_inst_ack_0 : boolean;
  signal type_cast_1540_inst_req_1 : boolean;
  signal type_cast_1540_inst_ack_1 : boolean;
  signal if_stmt_1553_branch_req_0 : boolean;
  signal if_stmt_1553_branch_ack_1 : boolean;
  signal if_stmt_1553_branch_ack_0 : boolean;
  signal type_cast_1581_inst_req_0 : boolean;
  signal type_cast_1581_inst_ack_0 : boolean;
  signal type_cast_1581_inst_req_1 : boolean;
  signal type_cast_1581_inst_ack_1 : boolean;
  signal type_cast_1597_inst_req_0 : boolean;
  signal type_cast_1597_inst_ack_0 : boolean;
  signal type_cast_1597_inst_req_1 : boolean;
  signal type_cast_1597_inst_ack_1 : boolean;
  signal if_stmt_1604_branch_req_0 : boolean;
  signal if_stmt_1604_branch_ack_1 : boolean;
  signal if_stmt_1604_branch_ack_0 : boolean;
  signal WPIPE_Block0_done_1640_inst_req_0 : boolean;
  signal WPIPE_Block0_done_1640_inst_ack_0 : boolean;
  signal WPIPE_Block0_done_1640_inst_req_1 : boolean;
  signal WPIPE_Block0_done_1640_inst_ack_1 : boolean;
  signal phi_stmt_1423_req_0 : boolean;
  signal phi_stmt_1402_req_0 : boolean;
  signal phi_stmt_1409_req_0 : boolean;
  signal phi_stmt_1416_req_0 : boolean;
  signal type_cast_1429_inst_req_0 : boolean;
  signal type_cast_1429_inst_ack_0 : boolean;
  signal type_cast_1429_inst_req_1 : boolean;
  signal type_cast_1429_inst_ack_1 : boolean;
  signal phi_stmt_1423_req_1 : boolean;
  signal type_cast_1408_inst_req_0 : boolean;
  signal type_cast_1408_inst_ack_0 : boolean;
  signal type_cast_1408_inst_req_1 : boolean;
  signal type_cast_1408_inst_ack_1 : boolean;
  signal phi_stmt_1402_req_1 : boolean;
  signal type_cast_1415_inst_req_0 : boolean;
  signal type_cast_1415_inst_ack_0 : boolean;
  signal type_cast_1415_inst_req_1 : boolean;
  signal type_cast_1415_inst_ack_1 : boolean;
  signal phi_stmt_1409_req_1 : boolean;
  signal type_cast_1422_inst_req_0 : boolean;
  signal type_cast_1422_inst_ack_0 : boolean;
  signal type_cast_1422_inst_req_1 : boolean;
  signal type_cast_1422_inst_ack_1 : boolean;
  signal phi_stmt_1416_req_1 : boolean;
  signal phi_stmt_1402_ack_0 : boolean;
  signal phi_stmt_1409_ack_0 : boolean;
  signal phi_stmt_1416_ack_0 : boolean;
  signal phi_stmt_1423_ack_0 : boolean;
  signal phi_stmt_1611_req_1 : boolean;
  signal type_cast_1623_inst_req_0 : boolean;
  signal type_cast_1623_inst_ack_0 : boolean;
  signal type_cast_1623_inst_req_1 : boolean;
  signal type_cast_1623_inst_ack_1 : boolean;
  signal phi_stmt_1618_req_1 : boolean;
  signal type_cast_1629_inst_req_0 : boolean;
  signal type_cast_1629_inst_ack_0 : boolean;
  signal type_cast_1629_inst_req_1 : boolean;
  signal type_cast_1629_inst_ack_1 : boolean;
  signal phi_stmt_1624_req_1 : boolean;
  signal type_cast_1614_inst_req_0 : boolean;
  signal type_cast_1614_inst_ack_0 : boolean;
  signal type_cast_1614_inst_req_1 : boolean;
  signal type_cast_1614_inst_ack_1 : boolean;
  signal phi_stmt_1611_req_0 : boolean;
  signal type_cast_1621_inst_req_0 : boolean;
  signal type_cast_1621_inst_ack_0 : boolean;
  signal type_cast_1621_inst_req_1 : boolean;
  signal type_cast_1621_inst_ack_1 : boolean;
  signal phi_stmt_1618_req_0 : boolean;
  signal type_cast_1627_inst_req_0 : boolean;
  signal type_cast_1627_inst_ack_0 : boolean;
  signal type_cast_1627_inst_req_1 : boolean;
  signal type_cast_1627_inst_ack_1 : boolean;
  signal phi_stmt_1624_req_0 : boolean;
  signal phi_stmt_1611_ack_0 : boolean;
  signal phi_stmt_1618_ack_0 : boolean;
  signal phi_stmt_1624_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeA_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeA_CP_3054_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeA_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_3054_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeA_CP_3054_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_3054_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeA_CP_3054: Block -- control-path 
    signal convTransposeA_CP_3054_elements: BooleanArray(125 downto 0);
    -- 
  begin -- 
    convTransposeA_CP_3054_elements(0) <= convTransposeA_CP_3054_start;
    convTransposeA_CP_3054_symbol <= convTransposeA_CP_3054_elements(78);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/type_cast_1326_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/type_cast_1339_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/type_cast_1326_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/type_cast_1339_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/type_cast_1339_Update/cr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1293/$entry
      -- CP-element group 0: 	 branch_block_stmt_1293/branch_block_stmt_1293__entry__
      -- CP-element group 0: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354__entry__
      -- CP-element group 0: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/$entry
      -- CP-element group 0: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1295_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1295_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1295_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/type_cast_1326_update_start_
      -- 
    cr_3247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(0), ack => type_cast_1326_inst_req_1); -- 
    cr_3275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(0), ack => type_cast_1339_inst_req_1); -- 
    rr_3102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(0), ack => RPIPE_Block0_start_1295_inst_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	125 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	84 
    -- CP-element group 1: 	85 
    -- CP-element group 1: 	87 
    -- CP-element group 1: 	88 
    -- CP-element group 1: 	90 
    -- CP-element group 1: 	91 
    -- CP-element group 1: 	93 
    -- CP-element group 1: 	94 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_1293/merge_stmt_1610__exit__
      -- CP-element group 1: 	 branch_block_stmt_1293/assign_stmt_1636__entry__
      -- CP-element group 1: 	 branch_block_stmt_1293/assign_stmt_1636__exit__
      -- CP-element group 1: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_1293/assign_stmt_1636/$entry
      -- CP-element group 1: 	 branch_block_stmt_1293/assign_stmt_1636/$exit
      -- CP-element group 1: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1423/$entry
      -- CP-element group 1: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1429/$entry
      -- CP-element group 1: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1429/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1429/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1429/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1429/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1429/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1402/$entry
      -- CP-element group 1: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1402/phi_stmt_1402_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1402/phi_stmt_1402_sources/type_cast_1408/$entry
      -- CP-element group 1: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1402/phi_stmt_1402_sources/type_cast_1408/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1402/phi_stmt_1402_sources/type_cast_1408/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1402/phi_stmt_1402_sources/type_cast_1408/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1402/phi_stmt_1402_sources/type_cast_1408/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1402/phi_stmt_1402_sources/type_cast_1408/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1409/$entry
      -- CP-element group 1: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1409/phi_stmt_1409_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1409/phi_stmt_1409_sources/type_cast_1415/$entry
      -- CP-element group 1: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1409/phi_stmt_1409_sources/type_cast_1415/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1409/phi_stmt_1409_sources/type_cast_1415/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1409/phi_stmt_1409_sources/type_cast_1415/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1409/phi_stmt_1409_sources/type_cast_1415/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1409/phi_stmt_1409_sources/type_cast_1415/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1416/$entry
      -- CP-element group 1: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1416/phi_stmt_1416_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1416/phi_stmt_1416_sources/type_cast_1422/$entry
      -- CP-element group 1: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1416/phi_stmt_1416_sources/type_cast_1422/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1416/phi_stmt_1416_sources/type_cast_1422/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1416/phi_stmt_1416_sources/type_cast_1422/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1416/phi_stmt_1416_sources/type_cast_1422/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1416/phi_stmt_1416_sources/type_cast_1422/SplitProtocol/Update/cr
      -- 
    rr_3788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(1), ack => type_cast_1429_inst_req_0); -- 
    cr_3793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(1), ack => type_cast_1429_inst_req_1); -- 
    rr_3811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(1), ack => type_cast_1408_inst_req_0); -- 
    cr_3816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(1), ack => type_cast_1408_inst_req_1); -- 
    rr_3834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(1), ack => type_cast_1415_inst_req_0); -- 
    cr_3839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(1), ack => type_cast_1415_inst_req_1); -- 
    rr_3857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(1), ack => type_cast_1422_inst_req_0); -- 
    cr_3862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(1), ack => type_cast_1422_inst_req_1); -- 
    convTransposeA_CP_3054_elements(1) <= convTransposeA_CP_3054_elements(125);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1295_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1295_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1295_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1295_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1295_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1295_Update/cr
      -- 
    ra_3103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1295_inst_ack_0, ack => convTransposeA_CP_3054_elements(2)); -- 
    cr_3107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(2), ack => RPIPE_Block0_start_1295_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1295_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1295_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1295_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1298_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1298_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1298_Sample/rr
      -- 
    ca_3108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1295_inst_ack_1, ack => convTransposeA_CP_3054_elements(3)); -- 
    rr_3116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(3), ack => RPIPE_Block0_start_1298_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1298_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1298_update_start_
      -- CP-element group 4: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1298_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1298_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1298_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1298_Update/cr
      -- 
    ra_3117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1298_inst_ack_0, ack => convTransposeA_CP_3054_elements(4)); -- 
    cr_3121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(4), ack => RPIPE_Block0_start_1298_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1298_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1298_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1298_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1301_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1301_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1301_Sample/rr
      -- 
    ca_3122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1298_inst_ack_1, ack => convTransposeA_CP_3054_elements(5)); -- 
    rr_3130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(5), ack => RPIPE_Block0_start_1301_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1301_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1301_update_start_
      -- CP-element group 6: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1301_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1301_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1301_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1301_Update/cr
      -- 
    ra_3131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1301_inst_ack_0, ack => convTransposeA_CP_3054_elements(6)); -- 
    cr_3135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(6), ack => RPIPE_Block0_start_1301_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1301_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1301_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1301_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1304_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1304_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1304_Sample/rr
      -- 
    ca_3136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1301_inst_ack_1, ack => convTransposeA_CP_3054_elements(7)); -- 
    rr_3144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(7), ack => RPIPE_Block0_start_1304_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1304_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1304_update_start_
      -- CP-element group 8: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1304_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1304_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1304_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1304_Update/cr
      -- 
    ra_3145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1304_inst_ack_0, ack => convTransposeA_CP_3054_elements(8)); -- 
    cr_3149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(8), ack => RPIPE_Block0_start_1304_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1304_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1304_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1304_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1307_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1307_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1307_Sample/rr
      -- 
    ca_3150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1304_inst_ack_1, ack => convTransposeA_CP_3054_elements(9)); -- 
    rr_3158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(9), ack => RPIPE_Block0_start_1307_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1307_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1307_update_start_
      -- CP-element group 10: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1307_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1307_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1307_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1307_Update/cr
      -- 
    ra_3159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1307_inst_ack_0, ack => convTransposeA_CP_3054_elements(10)); -- 
    cr_3163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(10), ack => RPIPE_Block0_start_1307_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1307_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1307_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1307_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1310_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1310_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1310_Sample/rr
      -- 
    ca_3164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1307_inst_ack_1, ack => convTransposeA_CP_3054_elements(11)); -- 
    rr_3172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(11), ack => RPIPE_Block0_start_1310_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1310_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1310_update_start_
      -- CP-element group 12: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1310_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1310_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1310_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1310_Update/cr
      -- 
    ra_3173_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1310_inst_ack_0, ack => convTransposeA_CP_3054_elements(12)); -- 
    cr_3177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(12), ack => RPIPE_Block0_start_1310_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1310_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1310_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1310_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1313_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1313_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1313_Sample/rr
      -- 
    ca_3178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1310_inst_ack_1, ack => convTransposeA_CP_3054_elements(13)); -- 
    rr_3186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(13), ack => RPIPE_Block0_start_1313_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1313_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1313_update_start_
      -- CP-element group 14: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1313_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1313_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1313_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1313_Update/cr
      -- 
    ra_3187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1313_inst_ack_0, ack => convTransposeA_CP_3054_elements(14)); -- 
    cr_3191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(14), ack => RPIPE_Block0_start_1313_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1313_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1313_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1313_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1316_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1316_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1316_Sample/rr
      -- 
    ca_3192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1313_inst_ack_1, ack => convTransposeA_CP_3054_elements(15)); -- 
    rr_3200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(15), ack => RPIPE_Block0_start_1316_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1316_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1316_update_start_
      -- CP-element group 16: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1316_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1316_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1316_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1316_Update/cr
      -- 
    ra_3201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1316_inst_ack_0, ack => convTransposeA_CP_3054_elements(16)); -- 
    cr_3205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(16), ack => RPIPE_Block0_start_1316_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1316_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1316_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1316_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1319_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1319_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1319_Sample/rr
      -- 
    ca_3206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1316_inst_ack_1, ack => convTransposeA_CP_3054_elements(17)); -- 
    rr_3214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(17), ack => RPIPE_Block0_start_1319_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1319_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1319_update_start_
      -- CP-element group 18: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1319_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1319_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1319_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1319_Update/cr
      -- 
    ra_3215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1319_inst_ack_0, ack => convTransposeA_CP_3054_elements(18)); -- 
    cr_3219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(18), ack => RPIPE_Block0_start_1319_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1319_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1319_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1319_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1322_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1322_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1322_Sample/rr
      -- 
    ca_3220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1319_inst_ack_1, ack => convTransposeA_CP_3054_elements(19)); -- 
    rr_3228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(19), ack => RPIPE_Block0_start_1322_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1322_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1322_update_start_
      -- CP-element group 20: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1322_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1322_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1322_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1322_Update/cr
      -- 
    ra_3229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1322_inst_ack_0, ack => convTransposeA_CP_3054_elements(20)); -- 
    cr_3233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(20), ack => RPIPE_Block0_start_1322_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1335_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1335_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1335_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1322_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1322_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1322_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/type_cast_1326_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/type_cast_1326_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/type_cast_1326_Sample/rr
      -- 
    ca_3234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1322_inst_ack_1, ack => convTransposeA_CP_3054_elements(21)); -- 
    rr_3242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(21), ack => type_cast_1326_inst_req_0); -- 
    rr_3256_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3256_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(21), ack => RPIPE_Block0_start_1335_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/type_cast_1326_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/type_cast_1326_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/type_cast_1326_Sample/ra
      -- 
    ra_3243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1326_inst_ack_0, ack => convTransposeA_CP_3054_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/type_cast_1326_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/type_cast_1326_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/type_cast_1326_update_completed_
      -- 
    ca_3248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1326_inst_ack_1, ack => convTransposeA_CP_3054_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1335_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1335_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1335_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1335_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1335_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1335_Update/cr
      -- 
    ra_3257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1335_inst_ack_0, ack => convTransposeA_CP_3054_elements(24)); -- 
    cr_3261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(24), ack => RPIPE_Block0_start_1335_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/type_cast_1339_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1335_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1347_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1347_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/type_cast_1339_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1335_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1347_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1335_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/type_cast_1339_sample_start_
      -- 
    ca_3262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1335_inst_ack_1, ack => convTransposeA_CP_3054_elements(25)); -- 
    rr_3270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(25), ack => type_cast_1339_inst_req_0); -- 
    rr_3284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(25), ack => RPIPE_Block0_start_1347_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/type_cast_1339_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/type_cast_1339_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/type_cast_1339_Sample/$exit
      -- 
    ra_3271_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1339_inst_ack_0, ack => convTransposeA_CP_3054_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/type_cast_1339_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/type_cast_1339_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/type_cast_1339_Update/ca
      -- 
    ca_3276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1339_inst_ack_1, ack => convTransposeA_CP_3054_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1347_Update/cr
      -- CP-element group 28: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1347_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1347_update_start_
      -- CP-element group 28: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1347_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1347_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1347_Sample/$exit
      -- 
    ra_3285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1347_inst_ack_0, ack => convTransposeA_CP_3054_elements(28)); -- 
    cr_3289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(28), ack => RPIPE_Block0_start_1347_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1347_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1350_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1350_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1350_Sample/rr
      -- CP-element group 29: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1347_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1347_Update/$exit
      -- 
    ca_3290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1347_inst_ack_1, ack => convTransposeA_CP_3054_elements(29)); -- 
    rr_3298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(29), ack => RPIPE_Block0_start_1350_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1350_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1350_update_start_
      -- CP-element group 30: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1350_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1350_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1350_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1350_Update/cr
      -- 
    ra_3299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1350_inst_ack_0, ack => convTransposeA_CP_3054_elements(30)); -- 
    cr_3303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(30), ack => RPIPE_Block0_start_1350_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1353_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1350_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1353_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1353_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1350_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1350_Update/ca
      -- 
    ca_3304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1350_inst_ack_1, ack => convTransposeA_CP_3054_elements(31)); -- 
    rr_3312_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3312_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(31), ack => RPIPE_Block0_start_1353_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1353_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1353_update_start_
      -- CP-element group 32: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1353_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1353_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1353_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1353_Update/cr
      -- 
    ra_3313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1353_inst_ack_0, ack => convTransposeA_CP_3054_elements(32)); -- 
    cr_3317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(32), ack => RPIPE_Block0_start_1353_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1353_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1353_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/RPIPE_Block0_start_1353_Update/ca
      -- 
    ca_3318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1353_inst_ack_1, ack => convTransposeA_CP_3054_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34: 	41 
    -- CP-element group 34: 	42 
    -- CP-element group 34:  members (28) 
      -- CP-element group 34: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1380_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1384_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1392_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1380_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1380_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1392_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1384_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1388_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1380_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1392_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1388_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1380_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1384_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1388_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1384_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1392_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1392_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1388_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1384_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1392_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1388_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1380_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1384_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/$entry
      -- CP-element group 34: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354__exit__
      -- CP-element group 34: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399__entry__
      -- CP-element group 34: 	 branch_block_stmt_1293/assign_stmt_1296_to_assign_stmt_1354/$exit
      -- CP-element group 34: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1388_Update/cr
      -- 
    rr_3329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(34), ack => type_cast_1380_inst_req_0); -- 
    cr_3376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(34), ack => type_cast_1392_inst_req_1); -- 
    cr_3334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(34), ack => type_cast_1380_inst_req_1); -- 
    rr_3343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(34), ack => type_cast_1384_inst_req_0); -- 
    rr_3371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(34), ack => type_cast_1392_inst_req_0); -- 
    rr_3357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(34), ack => type_cast_1388_inst_req_0); -- 
    cr_3348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(34), ack => type_cast_1384_inst_req_1); -- 
    cr_3362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(34), ack => type_cast_1388_inst_req_1); -- 
    convTransposeA_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3054_elements(23) & convTransposeA_CP_3054_elements(27) & convTransposeA_CP_3054_elements(33);
      gj_convTransposeA_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3054_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1380_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1380_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1380_Sample/$exit
      -- 
    ra_3330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1380_inst_ack_0, ack => convTransposeA_CP_3054_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	43 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1380_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1380_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1380_update_completed_
      -- 
    ca_3335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1380_inst_ack_1, ack => convTransposeA_CP_3054_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1384_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1384_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1384_sample_completed_
      -- 
    ra_3344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1384_inst_ack_0, ack => convTransposeA_CP_3054_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	43 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1384_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1384_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1384_Update/$exit
      -- 
    ca_3349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1384_inst_ack_1, ack => convTransposeA_CP_3054_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1388_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1388_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1388_Sample/ra
      -- 
    ra_3358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1388_inst_ack_0, ack => convTransposeA_CP_3054_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	43 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1388_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1388_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1388_Update/$exit
      -- 
    ca_3363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1388_inst_ack_1, ack => convTransposeA_CP_3054_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	34 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1392_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1392_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1392_Sample/ra
      -- 
    ra_3372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1392_inst_ack_0, ack => convTransposeA_CP_3054_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	34 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1392_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1392_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/type_cast_1392_Update/$exit
      -- 
    ca_3377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1392_inst_ack_1, ack => convTransposeA_CP_3054_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  place  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	36 
    -- CP-element group 43: 	38 
    -- CP-element group 43: 	40 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	79 
    -- CP-element group 43: 	80 
    -- CP-element group 43: 	81 
    -- CP-element group 43: 	82 
    -- CP-element group 43:  members (12) 
      -- CP-element group 43: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399/$exit
      -- CP-element group 43: 	 branch_block_stmt_1293/assign_stmt_1361_to_assign_stmt_1399__exit__
      -- CP-element group 43: 	 branch_block_stmt_1293/entry_whilex_xbody
      -- CP-element group 43: 	 branch_block_stmt_1293/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 43: 	 branch_block_stmt_1293/entry_whilex_xbody_PhiReq/phi_stmt_1423/$entry
      -- CP-element group 43: 	 branch_block_stmt_1293/entry_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1293/entry_whilex_xbody_PhiReq/phi_stmt_1402/$entry
      -- CP-element group 43: 	 branch_block_stmt_1293/entry_whilex_xbody_PhiReq/phi_stmt_1402/phi_stmt_1402_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1293/entry_whilex_xbody_PhiReq/phi_stmt_1409/$entry
      -- CP-element group 43: 	 branch_block_stmt_1293/entry_whilex_xbody_PhiReq/phi_stmt_1409/phi_stmt_1409_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1293/entry_whilex_xbody_PhiReq/phi_stmt_1416/$entry
      -- CP-element group 43: 	 branch_block_stmt_1293/entry_whilex_xbody_PhiReq/phi_stmt_1416/phi_stmt_1416_sources/$entry
      -- 
    convTransposeA_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3054_elements(36) & convTransposeA_CP_3054_elements(38) & convTransposeA_CP_3054_elements(40) & convTransposeA_CP_3054_elements(42);
      gj_convTransposeA_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3054_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	102 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1464_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1464_Sample/ra
      -- CP-element group 44: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1464_sample_completed_
      -- 
    ra_3389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1464_inst_ack_0, ack => convTransposeA_CP_3054_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	102 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	58 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1464_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1464_Update/ca
      -- CP-element group 45: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1464_update_completed_
      -- 
    ca_3394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1464_inst_ack_1, ack => convTransposeA_CP_3054_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	102 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1468_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1468_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1468_Sample/ra
      -- 
    ra_3403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1468_inst_ack_0, ack => convTransposeA_CP_3054_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	102 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	58 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1468_Update/ca
      -- CP-element group 47: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1468_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1468_Update/$exit
      -- 
    ca_3408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1468_inst_ack_1, ack => convTransposeA_CP_3054_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	102 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1472_Sample/ra
      -- CP-element group 48: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1472_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1472_sample_completed_
      -- 
    ra_3417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1472_inst_ack_0, ack => convTransposeA_CP_3054_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	102 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1472_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1472_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1472_Update/ca
      -- 
    ca_3422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1472_inst_ack_1, ack => convTransposeA_CP_3054_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	102 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1502_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1502_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1502_Sample/ra
      -- 
    ra_3431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1502_inst_ack_0, ack => convTransposeA_CP_3054_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	102 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (16) 
      -- CP-element group 51: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1502_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1502_Update/ca
      -- CP-element group 51: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1508_index_resized_1
      -- CP-element group 51: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1508_index_scaled_1
      -- CP-element group 51: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1502_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1508_index_computed_1
      -- CP-element group 51: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1508_index_resize_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1508_index_resize_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1508_index_resize_1/index_resize_req
      -- CP-element group 51: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1508_index_resize_1/index_resize_ack
      -- CP-element group 51: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1508_index_scale_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1508_index_scale_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1508_index_scale_1/scale_rename_req
      -- CP-element group 51: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1508_index_scale_1/scale_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1508_final_index_sum_regn_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1508_final_index_sum_regn_Sample/req
      -- 
    ca_3436_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1502_inst_ack_1, ack => convTransposeA_CP_3054_elements(51)); -- 
    req_3461_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3461_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(51), ack => array_obj_ref_1508_index_offset_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	68 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1508_final_index_sum_regn_sample_complete
      -- CP-element group 52: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1508_final_index_sum_regn_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1508_final_index_sum_regn_Sample/ack
      -- 
    ack_3462_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1508_index_offset_ack_0, ack => convTransposeA_CP_3054_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	102 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (11) 
      -- CP-element group 53: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/addr_of_1509_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1508_root_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1508_offset_calculated
      -- CP-element group 53: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1508_final_index_sum_regn_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1508_final_index_sum_regn_Update/ack
      -- CP-element group 53: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1508_base_plus_offset/$entry
      -- CP-element group 53: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1508_base_plus_offset/$exit
      -- CP-element group 53: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1508_base_plus_offset/sum_rename_req
      -- CP-element group 53: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1508_base_plus_offset/sum_rename_ack
      -- CP-element group 53: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/addr_of_1509_request/$entry
      -- CP-element group 53: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/addr_of_1509_request/req
      -- 
    ack_3467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1508_index_offset_ack_1, ack => convTransposeA_CP_3054_elements(53)); -- 
    req_3476_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3476_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(53), ack => addr_of_1509_final_reg_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/addr_of_1509_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/addr_of_1509_request/$exit
      -- CP-element group 54: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/addr_of_1509_request/ack
      -- 
    ack_3477_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1509_final_reg_ack_0, ack => convTransposeA_CP_3054_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	102 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (24) 
      -- CP-element group 55: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/addr_of_1509_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/addr_of_1509_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/addr_of_1509_complete/ack
      -- CP-element group 55: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1513_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1513_base_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1513_word_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1513_root_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1513_base_address_resized
      -- CP-element group 55: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1513_base_addr_resize/$entry
      -- CP-element group 55: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1513_base_addr_resize/$exit
      -- CP-element group 55: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1513_base_addr_resize/base_resize_req
      -- CP-element group 55: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1513_base_addr_resize/base_resize_ack
      -- CP-element group 55: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1513_base_plus_offset/$entry
      -- CP-element group 55: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1513_base_plus_offset/$exit
      -- CP-element group 55: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1513_base_plus_offset/sum_rename_req
      -- CP-element group 55: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1513_base_plus_offset/sum_rename_ack
      -- CP-element group 55: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1513_word_addrgen/$entry
      -- CP-element group 55: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1513_word_addrgen/$exit
      -- CP-element group 55: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1513_word_addrgen/root_register_req
      -- CP-element group 55: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1513_word_addrgen/root_register_ack
      -- CP-element group 55: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1513_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1513_Sample/word_access_start/$entry
      -- CP-element group 55: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1513_Sample/word_access_start/word_0/$entry
      -- CP-element group 55: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1513_Sample/word_access_start/word_0/rr
      -- 
    ack_3482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1509_final_reg_ack_1, ack => convTransposeA_CP_3054_elements(55)); -- 
    rr_3515_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3515_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(55), ack => ptr_deref_1513_load_0_req_0); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (5) 
      -- CP-element group 56: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1513_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1513_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1513_Sample/word_access_start/$exit
      -- CP-element group 56: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1513_Sample/word_access_start/word_0/$exit
      -- CP-element group 56: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1513_Sample/word_access_start/word_0/ra
      -- 
    ra_3516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1513_load_0_ack_0, ack => convTransposeA_CP_3054_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	102 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (9) 
      -- CP-element group 57: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1513_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1513_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1513_Update/word_access_complete/$exit
      -- CP-element group 57: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1513_Update/word_access_complete/word_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1513_Update/word_access_complete/word_0/ca
      -- CP-element group 57: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1513_Update/ptr_deref_1513_Merge/$entry
      -- CP-element group 57: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1513_Update/ptr_deref_1513_Merge/$exit
      -- CP-element group 57: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1513_Update/ptr_deref_1513_Merge/merge_req
      -- CP-element group 57: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1513_Update/ptr_deref_1513_Merge/merge_ack
      -- 
    ca_3527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1513_load_0_ack_1, ack => convTransposeA_CP_3054_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	45 
    -- CP-element group 58: 	47 
    -- CP-element group 58: 	49 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (13) 
      -- CP-element group 58: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1531_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1531_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1531_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1531_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1531_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1531_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1531_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1531_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1531_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1531_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1531_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1531_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1531_final_index_sum_regn_Sample/req
      -- 
    req_3557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(58), ack => array_obj_ref_1531_index_offset_req_0); -- 
    convTransposeA_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3054_elements(45) & convTransposeA_CP_3054_elements(47) & convTransposeA_CP_3054_elements(49);
      gj_convTransposeA_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3054_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	68 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1531_final_index_sum_regn_sample_complete
      -- CP-element group 59: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1531_final_index_sum_regn_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1531_final_index_sum_regn_Sample/ack
      -- 
    ack_3558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1531_index_offset_ack_0, ack => convTransposeA_CP_3054_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	102 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (11) 
      -- CP-element group 60: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/addr_of_1532_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1531_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1531_offset_calculated
      -- CP-element group 60: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1531_final_index_sum_regn_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1531_final_index_sum_regn_Update/ack
      -- CP-element group 60: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1531_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1531_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1531_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1531_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/addr_of_1532_request/$entry
      -- CP-element group 60: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/addr_of_1532_request/req
      -- 
    ack_3563_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1531_index_offset_ack_1, ack => convTransposeA_CP_3054_elements(60)); -- 
    req_3572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(60), ack => addr_of_1532_final_reg_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/addr_of_1532_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/addr_of_1532_request/$exit
      -- CP-element group 61: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/addr_of_1532_request/ack
      -- 
    ack_3573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1532_final_reg_ack_0, ack => convTransposeA_CP_3054_elements(61)); -- 
    -- CP-element group 62:  fork  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	102 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (19) 
      -- CP-element group 62: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/addr_of_1532_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/addr_of_1532_complete/$exit
      -- CP-element group 62: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/addr_of_1532_complete/ack
      -- CP-element group 62: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1535_base_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1535_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1535_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1535_base_address_resized
      -- CP-element group 62: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1535_base_addr_resize/$entry
      -- CP-element group 62: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1535_base_addr_resize/$exit
      -- CP-element group 62: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1535_base_addr_resize/base_resize_req
      -- CP-element group 62: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1535_base_addr_resize/base_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1535_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1535_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1535_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1535_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1535_word_addrgen/$entry
      -- CP-element group 62: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1535_word_addrgen/$exit
      -- CP-element group 62: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1535_word_addrgen/root_register_req
      -- CP-element group 62: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1535_word_addrgen/root_register_ack
      -- 
    ack_3578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1532_final_reg_ack_1, ack => convTransposeA_CP_3054_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1535_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1535_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1535_Sample/ptr_deref_1535_Split/$entry
      -- CP-element group 63: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1535_Sample/ptr_deref_1535_Split/$exit
      -- CP-element group 63: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1535_Sample/ptr_deref_1535_Split/split_req
      -- CP-element group 63: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1535_Sample/ptr_deref_1535_Split/split_ack
      -- CP-element group 63: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1535_Sample/word_access_start/$entry
      -- CP-element group 63: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1535_Sample/word_access_start/word_0/$entry
      -- CP-element group 63: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1535_Sample/word_access_start/word_0/rr
      -- 
    rr_3616_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3616_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(63), ack => ptr_deref_1535_store_0_req_0); -- 
    convTransposeA_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3054_elements(57) & convTransposeA_CP_3054_elements(62);
      gj_convTransposeA_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3054_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1535_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1535_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1535_Sample/word_access_start/$exit
      -- CP-element group 64: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1535_Sample/word_access_start/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1535_Sample/word_access_start/word_0/ra
      -- 
    ra_3617_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1535_store_0_ack_0, ack => convTransposeA_CP_3054_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	102 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	68 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1535_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1535_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1535_Update/word_access_complete/$exit
      -- CP-element group 65: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1535_Update/word_access_complete/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1535_Update/word_access_complete/word_0/ca
      -- 
    ca_3628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1535_store_0_ack_1, ack => convTransposeA_CP_3054_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	102 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1540_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1540_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1540_Sample/ra
      -- 
    ra_3637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1540_inst_ack_0, ack => convTransposeA_CP_3054_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	102 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1540_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1540_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1540_Update/ca
      -- 
    ca_3642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1540_inst_ack_1, ack => convTransposeA_CP_3054_elements(67)); -- 
    -- CP-element group 68:  branch  join  transition  place  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	52 
    -- CP-element group 68: 	59 
    -- CP-element group 68: 	65 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (10) 
      -- CP-element group 68: 	 branch_block_stmt_1293/R_cmp_1554_place
      -- CP-element group 68: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/$exit
      -- CP-element group 68: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552__exit__
      -- CP-element group 68: 	 branch_block_stmt_1293/if_stmt_1553__entry__
      -- CP-element group 68: 	 branch_block_stmt_1293/if_stmt_1553_dead_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1293/if_stmt_1553_eval_test/$entry
      -- CP-element group 68: 	 branch_block_stmt_1293/if_stmt_1553_eval_test/$exit
      -- CP-element group 68: 	 branch_block_stmt_1293/if_stmt_1553_eval_test/branch_req
      -- CP-element group 68: 	 branch_block_stmt_1293/if_stmt_1553_if_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1293/if_stmt_1553_else_link/$entry
      -- 
    branch_req_3650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(68), ack => if_stmt_1553_branch_req_0); -- 
    convTransposeA_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3054_elements(52) & convTransposeA_CP_3054_elements(59) & convTransposeA_CP_3054_elements(65) & convTransposeA_CP_3054_elements(67);
      gj_convTransposeA_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3054_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	111 
    -- CP-element group 69: 	112 
    -- CP-element group 69: 	114 
    -- CP-element group 69: 	115 
    -- CP-element group 69: 	117 
    -- CP-element group 69: 	118 
    -- CP-element group 69:  members (40) 
      -- CP-element group 69: 	 branch_block_stmt_1293/merge_stmt_1559__exit__
      -- CP-element group 69: 	 branch_block_stmt_1293/assign_stmt_1565__entry__
      -- CP-element group 69: 	 branch_block_stmt_1293/assign_stmt_1565__exit__
      -- CP-element group 69: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123
      -- CP-element group 69: 	 branch_block_stmt_1293/if_stmt_1553_if_link/$exit
      -- CP-element group 69: 	 branch_block_stmt_1293/if_stmt_1553_if_link/if_choice_transition
      -- CP-element group 69: 	 branch_block_stmt_1293/whilex_xbody_ifx_xthen
      -- CP-element group 69: 	 branch_block_stmt_1293/assign_stmt_1565/$entry
      -- CP-element group 69: 	 branch_block_stmt_1293/assign_stmt_1565/$exit
      -- CP-element group 69: 	 branch_block_stmt_1293/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1293/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 69: 	 branch_block_stmt_1293/merge_stmt_1559_PhiReqMerge
      -- CP-element group 69: 	 branch_block_stmt_1293/merge_stmt_1559_PhiAck/$entry
      -- CP-element group 69: 	 branch_block_stmt_1293/merge_stmt_1559_PhiAck/$exit
      -- CP-element group 69: 	 branch_block_stmt_1293/merge_stmt_1559_PhiAck/dummy
      -- CP-element group 69: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1611/$entry
      -- CP-element group 69: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1611/phi_stmt_1611_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1611/phi_stmt_1611_sources/type_cast_1614/$entry
      -- CP-element group 69: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1611/phi_stmt_1611_sources/type_cast_1614/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1611/phi_stmt_1611_sources/type_cast_1614/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1611/phi_stmt_1611_sources/type_cast_1614/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1611/phi_stmt_1611_sources/type_cast_1614/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1611/phi_stmt_1611_sources/type_cast_1614/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1618/$entry
      -- CP-element group 69: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/type_cast_1621/$entry
      -- CP-element group 69: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/type_cast_1621/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/type_cast_1621/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/type_cast_1621/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/type_cast_1621/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/type_cast_1621/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1624/$entry
      -- CP-element group 69: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1627/$entry
      -- CP-element group 69: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1627/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1627/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1627/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1627/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1627/SplitProtocol/Update/cr
      -- 
    if_choice_transition_3655_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1553_branch_ack_1, ack => convTransposeA_CP_3054_elements(69)); -- 
    rr_3972_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3972_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(69), ack => type_cast_1614_inst_req_0); -- 
    cr_3977_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3977_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(69), ack => type_cast_1614_inst_req_1); -- 
    rr_3995_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3995_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(69), ack => type_cast_1621_inst_req_0); -- 
    cr_4000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(69), ack => type_cast_1621_inst_req_1); -- 
    rr_4018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(69), ack => type_cast_1627_inst_req_0); -- 
    cr_4023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(69), ack => type_cast_1627_inst_req_1); -- 
    -- CP-element group 70:  fork  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70: 	74 
    -- CP-element group 70:  members (21) 
      -- CP-element group 70: 	 branch_block_stmt_1293/merge_stmt_1567__exit__
      -- CP-element group 70: 	 branch_block_stmt_1293/assign_stmt_1573_to_assign_stmt_1603__entry__
      -- CP-element group 70: 	 branch_block_stmt_1293/if_stmt_1553_else_link/$exit
      -- CP-element group 70: 	 branch_block_stmt_1293/if_stmt_1553_else_link/else_choice_transition
      -- CP-element group 70: 	 branch_block_stmt_1293/whilex_xbody_ifx_xelse
      -- CP-element group 70: 	 branch_block_stmt_1293/assign_stmt_1573_to_assign_stmt_1603/$entry
      -- CP-element group 70: 	 branch_block_stmt_1293/assign_stmt_1573_to_assign_stmt_1603/type_cast_1581_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_1293/assign_stmt_1573_to_assign_stmt_1603/type_cast_1581_update_start_
      -- CP-element group 70: 	 branch_block_stmt_1293/assign_stmt_1573_to_assign_stmt_1603/type_cast_1581_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_1293/assign_stmt_1573_to_assign_stmt_1603/type_cast_1581_Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_1293/assign_stmt_1573_to_assign_stmt_1603/type_cast_1581_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1293/assign_stmt_1573_to_assign_stmt_1603/type_cast_1581_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_1293/assign_stmt_1573_to_assign_stmt_1603/type_cast_1597_update_start_
      -- CP-element group 70: 	 branch_block_stmt_1293/assign_stmt_1573_to_assign_stmt_1603/type_cast_1597_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1293/assign_stmt_1573_to_assign_stmt_1603/type_cast_1597_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_1293/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_1293/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 70: 	 branch_block_stmt_1293/merge_stmt_1567_PhiReqMerge
      -- CP-element group 70: 	 branch_block_stmt_1293/merge_stmt_1567_PhiAck/$entry
      -- CP-element group 70: 	 branch_block_stmt_1293/merge_stmt_1567_PhiAck/$exit
      -- CP-element group 70: 	 branch_block_stmt_1293/merge_stmt_1567_PhiAck/dummy
      -- 
    else_choice_transition_3659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1553_branch_ack_0, ack => convTransposeA_CP_3054_elements(70)); -- 
    rr_3675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(70), ack => type_cast_1581_inst_req_0); -- 
    cr_3680_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3680_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(70), ack => type_cast_1581_inst_req_1); -- 
    cr_3694_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3694_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(70), ack => type_cast_1597_inst_req_1); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_1293/assign_stmt_1573_to_assign_stmt_1603/type_cast_1581_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_1293/assign_stmt_1573_to_assign_stmt_1603/type_cast_1581_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_1293/assign_stmt_1573_to_assign_stmt_1603/type_cast_1581_Sample/ra
      -- 
    ra_3676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1581_inst_ack_0, ack => convTransposeA_CP_3054_elements(71)); -- 
    -- CP-element group 72:  transition  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (6) 
      -- CP-element group 72: 	 branch_block_stmt_1293/assign_stmt_1573_to_assign_stmt_1603/type_cast_1581_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_1293/assign_stmt_1573_to_assign_stmt_1603/type_cast_1581_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_1293/assign_stmt_1573_to_assign_stmt_1603/type_cast_1581_Update/ca
      -- CP-element group 72: 	 branch_block_stmt_1293/assign_stmt_1573_to_assign_stmt_1603/type_cast_1597_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_1293/assign_stmt_1573_to_assign_stmt_1603/type_cast_1597_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_1293/assign_stmt_1573_to_assign_stmt_1603/type_cast_1597_Sample/rr
      -- 
    ca_3681_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1581_inst_ack_1, ack => convTransposeA_CP_3054_elements(72)); -- 
    rr_3689_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3689_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(72), ack => type_cast_1597_inst_req_0); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1293/assign_stmt_1573_to_assign_stmt_1603/type_cast_1597_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_1293/assign_stmt_1573_to_assign_stmt_1603/type_cast_1597_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_1293/assign_stmt_1573_to_assign_stmt_1603/type_cast_1597_Sample/ra
      -- 
    ra_3690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1597_inst_ack_0, ack => convTransposeA_CP_3054_elements(73)); -- 
    -- CP-element group 74:  branch  transition  place  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	70 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (13) 
      -- CP-element group 74: 	 branch_block_stmt_1293/assign_stmt_1573_to_assign_stmt_1603__exit__
      -- CP-element group 74: 	 branch_block_stmt_1293/if_stmt_1604__entry__
      -- CP-element group 74: 	 branch_block_stmt_1293/assign_stmt_1573_to_assign_stmt_1603/$exit
      -- CP-element group 74: 	 branch_block_stmt_1293/assign_stmt_1573_to_assign_stmt_1603/type_cast_1597_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_1293/assign_stmt_1573_to_assign_stmt_1603/type_cast_1597_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_1293/assign_stmt_1573_to_assign_stmt_1603/type_cast_1597_Update/ca
      -- CP-element group 74: 	 branch_block_stmt_1293/if_stmt_1604_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1293/if_stmt_1604_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_1293/if_stmt_1604_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_1293/if_stmt_1604_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_1293/R_cmp112_1605_place
      -- CP-element group 74: 	 branch_block_stmt_1293/if_stmt_1604_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1293/if_stmt_1604_else_link/$entry
      -- 
    ca_3695_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1597_inst_ack_1, ack => convTransposeA_CP_3054_elements(74)); -- 
    branch_req_3703_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3703_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(74), ack => if_stmt_1604_branch_req_0); -- 
    -- CP-element group 75:  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (15) 
      -- CP-element group 75: 	 branch_block_stmt_1293/merge_stmt_1638__exit__
      -- CP-element group 75: 	 branch_block_stmt_1293/assign_stmt_1643__entry__
      -- CP-element group 75: 	 branch_block_stmt_1293/if_stmt_1604_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_1293/if_stmt_1604_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_1293/ifx_xelse_whilex_xend
      -- CP-element group 75: 	 branch_block_stmt_1293/assign_stmt_1643/$entry
      -- CP-element group 75: 	 branch_block_stmt_1293/assign_stmt_1643/WPIPE_Block0_done_1640_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_1293/assign_stmt_1643/WPIPE_Block0_done_1640_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_1293/assign_stmt_1643/WPIPE_Block0_done_1640_Sample/req
      -- CP-element group 75: 	 branch_block_stmt_1293/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_1293/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_1293/merge_stmt_1638_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_1293/merge_stmt_1638_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_1293/merge_stmt_1638_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_1293/merge_stmt_1638_PhiAck/dummy
      -- 
    if_choice_transition_3708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1604_branch_ack_1, ack => convTransposeA_CP_3054_elements(75)); -- 
    req_3728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(75), ack => WPIPE_Block0_done_1640_inst_req_0); -- 
    -- CP-element group 76:  fork  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	103 
    -- CP-element group 76: 	104 
    -- CP-element group 76: 	105 
    -- CP-element group 76: 	107 
    -- CP-element group 76: 	108 
    -- CP-element group 76:  members (22) 
      -- CP-element group 76: 	 branch_block_stmt_1293/if_stmt_1604_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_1293/if_stmt_1604_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123
      -- CP-element group 76: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1611/$entry
      -- CP-element group 76: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1611/phi_stmt_1611_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1618/$entry
      -- CP-element group 76: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/type_cast_1623/$entry
      -- CP-element group 76: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/type_cast_1623/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/type_cast_1623/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/type_cast_1623/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/type_cast_1623/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/type_cast_1623/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1624/$entry
      -- CP-element group 76: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1629/$entry
      -- CP-element group 76: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1629/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1629/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1629/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1629/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1629/SplitProtocol/Update/cr
      -- 
    else_choice_transition_3712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1604_branch_ack_0, ack => convTransposeA_CP_3054_elements(76)); -- 
    rr_3923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(76), ack => type_cast_1623_inst_req_0); -- 
    cr_3928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(76), ack => type_cast_1623_inst_req_1); -- 
    rr_3946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(76), ack => type_cast_1629_inst_req_0); -- 
    cr_3951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(76), ack => type_cast_1629_inst_req_1); -- 
    -- CP-element group 77:  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (6) 
      -- CP-element group 77: 	 branch_block_stmt_1293/assign_stmt_1643/WPIPE_Block0_done_1640_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_1293/assign_stmt_1643/WPIPE_Block0_done_1640_update_start_
      -- CP-element group 77: 	 branch_block_stmt_1293/assign_stmt_1643/WPIPE_Block0_done_1640_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_1293/assign_stmt_1643/WPIPE_Block0_done_1640_Sample/ack
      -- CP-element group 77: 	 branch_block_stmt_1293/assign_stmt_1643/WPIPE_Block0_done_1640_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1293/assign_stmt_1643/WPIPE_Block0_done_1640_Update/req
      -- 
    ack_3729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1640_inst_ack_0, ack => convTransposeA_CP_3054_elements(77)); -- 
    req_3733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(77), ack => WPIPE_Block0_done_1640_inst_req_1); -- 
    -- CP-element group 78:  transition  place  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (16) 
      -- CP-element group 78: 	 $exit
      -- CP-element group 78: 	 branch_block_stmt_1293/$exit
      -- CP-element group 78: 	 branch_block_stmt_1293/branch_block_stmt_1293__exit__
      -- CP-element group 78: 	 branch_block_stmt_1293/assign_stmt_1643__exit__
      -- CP-element group 78: 	 branch_block_stmt_1293/return__
      -- CP-element group 78: 	 branch_block_stmt_1293/merge_stmt_1645__exit__
      -- CP-element group 78: 	 branch_block_stmt_1293/assign_stmt_1643/$exit
      -- CP-element group 78: 	 branch_block_stmt_1293/assign_stmt_1643/WPIPE_Block0_done_1640_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_1293/assign_stmt_1643/WPIPE_Block0_done_1640_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_1293/assign_stmt_1643/WPIPE_Block0_done_1640_Update/ack
      -- CP-element group 78: 	 branch_block_stmt_1293/return___PhiReq/$entry
      -- CP-element group 78: 	 branch_block_stmt_1293/return___PhiReq/$exit
      -- CP-element group 78: 	 branch_block_stmt_1293/merge_stmt_1645_PhiReqMerge
      -- CP-element group 78: 	 branch_block_stmt_1293/merge_stmt_1645_PhiAck/$entry
      -- CP-element group 78: 	 branch_block_stmt_1293/merge_stmt_1645_PhiAck/$exit
      -- CP-element group 78: 	 branch_block_stmt_1293/merge_stmt_1645_PhiAck/dummy
      -- 
    ack_3734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1640_inst_ack_1, ack => convTransposeA_CP_3054_elements(78)); -- 
    -- CP-element group 79:  transition  output  delay-element  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	43 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	83 
    -- CP-element group 79:  members (4) 
      -- CP-element group 79: 	 branch_block_stmt_1293/entry_whilex_xbody_PhiReq/phi_stmt_1423/$exit
      -- CP-element group 79: 	 branch_block_stmt_1293/entry_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/$exit
      -- CP-element group 79: 	 branch_block_stmt_1293/entry_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1427_konst_delay_trans
      -- CP-element group 79: 	 branch_block_stmt_1293/entry_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_req
      -- 
    phi_stmt_1423_req_3745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1423_req_3745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(79), ack => phi_stmt_1423_req_0); -- 
    -- Element group convTransposeA_CP_3054_elements(79) is a control-delay.
    cp_element_79_delay: control_delay_element  generic map(name => " 79_delay", delay_value => 1)  port map(req => convTransposeA_CP_3054_elements(43), ack => convTransposeA_CP_3054_elements(79), clk => clk, reset =>reset);
    -- CP-element group 80:  transition  output  delay-element  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	43 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	83 
    -- CP-element group 80:  members (4) 
      -- CP-element group 80: 	 branch_block_stmt_1293/entry_whilex_xbody_PhiReq/phi_stmt_1402/$exit
      -- CP-element group 80: 	 branch_block_stmt_1293/entry_whilex_xbody_PhiReq/phi_stmt_1402/phi_stmt_1402_sources/$exit
      -- CP-element group 80: 	 branch_block_stmt_1293/entry_whilex_xbody_PhiReq/phi_stmt_1402/phi_stmt_1402_sources/type_cast_1406_konst_delay_trans
      -- CP-element group 80: 	 branch_block_stmt_1293/entry_whilex_xbody_PhiReq/phi_stmt_1402/phi_stmt_1402_req
      -- 
    phi_stmt_1402_req_3753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1402_req_3753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(80), ack => phi_stmt_1402_req_0); -- 
    -- Element group convTransposeA_CP_3054_elements(80) is a control-delay.
    cp_element_80_delay: control_delay_element  generic map(name => " 80_delay", delay_value => 1)  port map(req => convTransposeA_CP_3054_elements(43), ack => convTransposeA_CP_3054_elements(80), clk => clk, reset =>reset);
    -- CP-element group 81:  transition  output  delay-element  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	43 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (4) 
      -- CP-element group 81: 	 branch_block_stmt_1293/entry_whilex_xbody_PhiReq/phi_stmt_1409/$exit
      -- CP-element group 81: 	 branch_block_stmt_1293/entry_whilex_xbody_PhiReq/phi_stmt_1409/phi_stmt_1409_sources/$exit
      -- CP-element group 81: 	 branch_block_stmt_1293/entry_whilex_xbody_PhiReq/phi_stmt_1409/phi_stmt_1409_sources/type_cast_1413_konst_delay_trans
      -- CP-element group 81: 	 branch_block_stmt_1293/entry_whilex_xbody_PhiReq/phi_stmt_1409/phi_stmt_1409_req
      -- 
    phi_stmt_1409_req_3761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1409_req_3761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(81), ack => phi_stmt_1409_req_0); -- 
    -- Element group convTransposeA_CP_3054_elements(81) is a control-delay.
    cp_element_81_delay: control_delay_element  generic map(name => " 81_delay", delay_value => 1)  port map(req => convTransposeA_CP_3054_elements(43), ack => convTransposeA_CP_3054_elements(81), clk => clk, reset =>reset);
    -- CP-element group 82:  transition  output  delay-element  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	43 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (4) 
      -- CP-element group 82: 	 branch_block_stmt_1293/entry_whilex_xbody_PhiReq/phi_stmt_1416/$exit
      -- CP-element group 82: 	 branch_block_stmt_1293/entry_whilex_xbody_PhiReq/phi_stmt_1416/phi_stmt_1416_sources/$exit
      -- CP-element group 82: 	 branch_block_stmt_1293/entry_whilex_xbody_PhiReq/phi_stmt_1416/phi_stmt_1416_sources/type_cast_1420_konst_delay_trans
      -- CP-element group 82: 	 branch_block_stmt_1293/entry_whilex_xbody_PhiReq/phi_stmt_1416/phi_stmt_1416_req
      -- 
    phi_stmt_1416_req_3769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1416_req_3769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(82), ack => phi_stmt_1416_req_0); -- 
    -- Element group convTransposeA_CP_3054_elements(82) is a control-delay.
    cp_element_82_delay: control_delay_element  generic map(name => " 82_delay", delay_value => 1)  port map(req => convTransposeA_CP_3054_elements(43), ack => convTransposeA_CP_3054_elements(82), clk => clk, reset =>reset);
    -- CP-element group 83:  join  transition  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	79 
    -- CP-element group 83: 	80 
    -- CP-element group 83: 	81 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	97 
    -- CP-element group 83:  members (1) 
      -- CP-element group 83: 	 branch_block_stmt_1293/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3054_elements(79) & convTransposeA_CP_3054_elements(80) & convTransposeA_CP_3054_elements(81) & convTransposeA_CP_3054_elements(82);
      gj_convTransposeA_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3054_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	1 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1429/SplitProtocol/Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1429/SplitProtocol/Sample/ra
      -- 
    ra_3789_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1429_inst_ack_0, ack => convTransposeA_CP_3054_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	1 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1429/SplitProtocol/Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1429/SplitProtocol/Update/ca
      -- 
    ca_3794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1429_inst_ack_1, ack => convTransposeA_CP_3054_elements(85)); -- 
    -- CP-element group 86:  join  transition  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	96 
    -- CP-element group 86:  members (5) 
      -- CP-element group 86: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1423/$exit
      -- CP-element group 86: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/$exit
      -- CP-element group 86: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1429/$exit
      -- CP-element group 86: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1429/SplitProtocol/$exit
      -- CP-element group 86: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_req
      -- 
    phi_stmt_1423_req_3795_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1423_req_3795_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(86), ack => phi_stmt_1423_req_1); -- 
    convTransposeA_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3054_elements(84) & convTransposeA_CP_3054_elements(85);
      gj_convTransposeA_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3054_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	1 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1402/phi_stmt_1402_sources/type_cast_1408/SplitProtocol/Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1402/phi_stmt_1402_sources/type_cast_1408/SplitProtocol/Sample/ra
      -- 
    ra_3812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1408_inst_ack_0, ack => convTransposeA_CP_3054_elements(87)); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	1 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1402/phi_stmt_1402_sources/type_cast_1408/SplitProtocol/Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1402/phi_stmt_1402_sources/type_cast_1408/SplitProtocol/Update/ca
      -- 
    ca_3817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1408_inst_ack_1, ack => convTransposeA_CP_3054_elements(88)); -- 
    -- CP-element group 89:  join  transition  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	96 
    -- CP-element group 89:  members (5) 
      -- CP-element group 89: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1402/$exit
      -- CP-element group 89: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1402/phi_stmt_1402_sources/$exit
      -- CP-element group 89: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1402/phi_stmt_1402_sources/type_cast_1408/$exit
      -- CP-element group 89: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1402/phi_stmt_1402_sources/type_cast_1408/SplitProtocol/$exit
      -- CP-element group 89: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1402/phi_stmt_1402_req
      -- 
    phi_stmt_1402_req_3818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1402_req_3818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(89), ack => phi_stmt_1402_req_1); -- 
    convTransposeA_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3054_elements(87) & convTransposeA_CP_3054_elements(88);
      gj_convTransposeA_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3054_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	1 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1409/phi_stmt_1409_sources/type_cast_1415/SplitProtocol/Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1409/phi_stmt_1409_sources/type_cast_1415/SplitProtocol/Sample/ra
      -- 
    ra_3835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1415_inst_ack_0, ack => convTransposeA_CP_3054_elements(90)); -- 
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	1 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1409/phi_stmt_1409_sources/type_cast_1415/SplitProtocol/Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1409/phi_stmt_1409_sources/type_cast_1415/SplitProtocol/Update/ca
      -- 
    ca_3840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1415_inst_ack_1, ack => convTransposeA_CP_3054_elements(91)); -- 
    -- CP-element group 92:  join  transition  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	96 
    -- CP-element group 92:  members (5) 
      -- CP-element group 92: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1409/$exit
      -- CP-element group 92: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1409/phi_stmt_1409_sources/$exit
      -- CP-element group 92: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1409/phi_stmt_1409_sources/type_cast_1415/$exit
      -- CP-element group 92: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1409/phi_stmt_1409_sources/type_cast_1415/SplitProtocol/$exit
      -- CP-element group 92: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1409/phi_stmt_1409_req
      -- 
    phi_stmt_1409_req_3841_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1409_req_3841_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(92), ack => phi_stmt_1409_req_1); -- 
    convTransposeA_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3054_elements(90) & convTransposeA_CP_3054_elements(91);
      gj_convTransposeA_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3054_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	1 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1416/phi_stmt_1416_sources/type_cast_1422/SplitProtocol/Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1416/phi_stmt_1416_sources/type_cast_1422/SplitProtocol/Sample/ra
      -- 
    ra_3858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1422_inst_ack_0, ack => convTransposeA_CP_3054_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	1 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1416/phi_stmt_1416_sources/type_cast_1422/SplitProtocol/Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1416/phi_stmt_1416_sources/type_cast_1422/SplitProtocol/Update/ca
      -- 
    ca_3863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1422_inst_ack_1, ack => convTransposeA_CP_3054_elements(94)); -- 
    -- CP-element group 95:  join  transition  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (5) 
      -- CP-element group 95: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1416/$exit
      -- CP-element group 95: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1416/phi_stmt_1416_sources/$exit
      -- CP-element group 95: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1416/phi_stmt_1416_sources/type_cast_1422/$exit
      -- CP-element group 95: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1416/phi_stmt_1416_sources/type_cast_1422/SplitProtocol/$exit
      -- CP-element group 95: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1416/phi_stmt_1416_req
      -- 
    phi_stmt_1416_req_3864_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1416_req_3864_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(95), ack => phi_stmt_1416_req_1); -- 
    convTransposeA_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3054_elements(93) & convTransposeA_CP_3054_elements(94);
      gj_convTransposeA_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3054_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  join  transition  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	86 
    -- CP-element group 96: 	89 
    -- CP-element group 96: 	92 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_1293/ifx_xend123_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3054_elements(86) & convTransposeA_CP_3054_elements(89) & convTransposeA_CP_3054_elements(92) & convTransposeA_CP_3054_elements(95);
      gj_convTransposeA_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3054_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  merge  fork  transition  place  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	83 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97: 	99 
    -- CP-element group 97: 	100 
    -- CP-element group 97: 	101 
    -- CP-element group 97:  members (2) 
      -- CP-element group 97: 	 branch_block_stmt_1293/merge_stmt_1401_PhiReqMerge
      -- CP-element group 97: 	 branch_block_stmt_1293/merge_stmt_1401_PhiAck/$entry
      -- 
    convTransposeA_CP_3054_elements(97) <= OrReduce(convTransposeA_CP_3054_elements(83) & convTransposeA_CP_3054_elements(96));
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	102 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_1293/merge_stmt_1401_PhiAck/phi_stmt_1402_ack
      -- 
    phi_stmt_1402_ack_3869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1402_ack_0, ack => convTransposeA_CP_3054_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	97 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	102 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_1293/merge_stmt_1401_PhiAck/phi_stmt_1409_ack
      -- 
    phi_stmt_1409_ack_3870_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1409_ack_0, ack => convTransposeA_CP_3054_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	97 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	102 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_1293/merge_stmt_1401_PhiAck/phi_stmt_1416_ack
      -- 
    phi_stmt_1416_ack_3871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1416_ack_0, ack => convTransposeA_CP_3054_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	97 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	102 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_1293/merge_stmt_1401_PhiAck/phi_stmt_1423_ack
      -- 
    phi_stmt_1423_ack_3872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1423_ack_0, ack => convTransposeA_CP_3054_elements(101)); -- 
    -- CP-element group 102:  join  fork  transition  place  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	98 
    -- CP-element group 102: 	99 
    -- CP-element group 102: 	100 
    -- CP-element group 102: 	101 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	44 
    -- CP-element group 102: 	45 
    -- CP-element group 102: 	46 
    -- CP-element group 102: 	47 
    -- CP-element group 102: 	48 
    -- CP-element group 102: 	49 
    -- CP-element group 102: 	50 
    -- CP-element group 102: 	51 
    -- CP-element group 102: 	53 
    -- CP-element group 102: 	55 
    -- CP-element group 102: 	57 
    -- CP-element group 102: 	60 
    -- CP-element group 102: 	62 
    -- CP-element group 102: 	65 
    -- CP-element group 102: 	66 
    -- CP-element group 102: 	67 
    -- CP-element group 102:  members (56) 
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1472_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1472_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1472_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1502_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1502_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1468_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/$entry
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1502_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1502_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1464_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/addr_of_1509_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1464_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1502_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1468_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1464_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1472_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1464_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1472_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1468_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1468_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1464_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1468_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1464_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1468_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1472_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1502_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1293/merge_stmt_1401__exit__
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552__entry__
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1508_final_index_sum_regn_update_start
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1508_final_index_sum_regn_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1508_final_index_sum_regn_Update/req
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/addr_of_1509_complete/$entry
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/addr_of_1509_complete/req
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1513_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1513_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1513_Update/word_access_complete/$entry
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1513_Update/word_access_complete/word_0/$entry
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1513_Update/word_access_complete/word_0/cr
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/addr_of_1532_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1531_final_index_sum_regn_update_start
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1531_final_index_sum_regn_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/array_obj_ref_1531_final_index_sum_regn_Update/req
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/addr_of_1532_complete/$entry
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/addr_of_1532_complete/req
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1535_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1535_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1535_Update/word_access_complete/$entry
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1535_Update/word_access_complete/word_0/$entry
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/ptr_deref_1535_Update/word_access_complete/word_0/cr
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1540_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1540_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1540_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1540_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1540_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1293/assign_stmt_1436_to_assign_stmt_1552/type_cast_1540_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1293/merge_stmt_1401_PhiAck/$exit
      -- 
    cr_3421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(102), ack => type_cast_1472_inst_req_1); -- 
    rr_3430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(102), ack => type_cast_1502_inst_req_0); -- 
    cr_3435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(102), ack => type_cast_1502_inst_req_1); -- 
    cr_3393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(102), ack => type_cast_1464_inst_req_1); -- 
    rr_3416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(102), ack => type_cast_1472_inst_req_0); -- 
    rr_3402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(102), ack => type_cast_1468_inst_req_0); -- 
    cr_3407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(102), ack => type_cast_1468_inst_req_1); -- 
    rr_3388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(102), ack => type_cast_1464_inst_req_0); -- 
    req_3466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(102), ack => array_obj_ref_1508_index_offset_req_1); -- 
    req_3481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(102), ack => addr_of_1509_final_reg_req_1); -- 
    cr_3526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(102), ack => ptr_deref_1513_load_0_req_1); -- 
    req_3562_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3562_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(102), ack => array_obj_ref_1531_index_offset_req_1); -- 
    req_3577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(102), ack => addr_of_1532_final_reg_req_1); -- 
    cr_3627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(102), ack => ptr_deref_1535_store_0_req_1); -- 
    rr_3636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(102), ack => type_cast_1540_inst_req_0); -- 
    cr_3641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(102), ack => type_cast_1540_inst_req_1); -- 
    convTransposeA_cp_element_group_102: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_102"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3054_elements(98) & convTransposeA_CP_3054_elements(99) & convTransposeA_CP_3054_elements(100) & convTransposeA_CP_3054_elements(101);
      gj_convTransposeA_cp_element_group_102 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3054_elements(102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 103:  transition  output  delay-element  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	76 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	110 
    -- CP-element group 103:  members (4) 
      -- CP-element group 103: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1611/$exit
      -- CP-element group 103: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1611/phi_stmt_1611_sources/$exit
      -- CP-element group 103: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1611/phi_stmt_1611_sources/type_cast_1617_konst_delay_trans
      -- CP-element group 103: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1611/phi_stmt_1611_req
      -- 
    phi_stmt_1611_req_3907_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1611_req_3907_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(103), ack => phi_stmt_1611_req_1); -- 
    -- Element group convTransposeA_CP_3054_elements(103) is a control-delay.
    cp_element_103_delay: control_delay_element  generic map(name => " 103_delay", delay_value => 1)  port map(req => convTransposeA_CP_3054_elements(76), ack => convTransposeA_CP_3054_elements(103), clk => clk, reset =>reset);
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	76 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	106 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/type_cast_1623/SplitProtocol/Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/type_cast_1623/SplitProtocol/Sample/ra
      -- 
    ra_3924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1623_inst_ack_0, ack => convTransposeA_CP_3054_elements(104)); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	76 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	106 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/type_cast_1623/SplitProtocol/Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/type_cast_1623/SplitProtocol/Update/ca
      -- 
    ca_3929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1623_inst_ack_1, ack => convTransposeA_CP_3054_elements(105)); -- 
    -- CP-element group 106:  join  transition  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	104 
    -- CP-element group 106: 	105 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	110 
    -- CP-element group 106:  members (5) 
      -- CP-element group 106: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1618/$exit
      -- CP-element group 106: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/$exit
      -- CP-element group 106: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/type_cast_1623/$exit
      -- CP-element group 106: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/type_cast_1623/SplitProtocol/$exit
      -- CP-element group 106: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1618/phi_stmt_1618_req
      -- 
    phi_stmt_1618_req_3930_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1618_req_3930_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(106), ack => phi_stmt_1618_req_1); -- 
    convTransposeA_cp_element_group_106: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_106"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3054_elements(104) & convTransposeA_CP_3054_elements(105);
      gj_convTransposeA_cp_element_group_106 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3054_elements(106), clk => clk, reset => reset); --
    end block;
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	76 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	109 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1629/SplitProtocol/Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1629/SplitProtocol/Sample/ra
      -- 
    ra_3947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1629_inst_ack_0, ack => convTransposeA_CP_3054_elements(107)); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	76 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (2) 
      -- CP-element group 108: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1629/SplitProtocol/Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1629/SplitProtocol/Update/ca
      -- 
    ca_3952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1629_inst_ack_1, ack => convTransposeA_CP_3054_elements(108)); -- 
    -- CP-element group 109:  join  transition  output  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	107 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109:  members (5) 
      -- CP-element group 109: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1624/$exit
      -- CP-element group 109: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/$exit
      -- CP-element group 109: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1629/$exit
      -- CP-element group 109: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1629/SplitProtocol/$exit
      -- CP-element group 109: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1624/phi_stmt_1624_req
      -- 
    phi_stmt_1624_req_3953_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1624_req_3953_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(109), ack => phi_stmt_1624_req_1); -- 
    convTransposeA_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3054_elements(107) & convTransposeA_CP_3054_elements(108);
      gj_convTransposeA_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3054_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  join  transition  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	103 
    -- CP-element group 110: 	106 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	121 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_1293/ifx_xelse_ifx_xend123_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3054_elements(103) & convTransposeA_CP_3054_elements(106) & convTransposeA_CP_3054_elements(109);
      gj_convTransposeA_cp_element_group_110 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3054_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	69 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	113 
    -- CP-element group 111:  members (2) 
      -- CP-element group 111: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1611/phi_stmt_1611_sources/type_cast_1614/SplitProtocol/Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1611/phi_stmt_1611_sources/type_cast_1614/SplitProtocol/Sample/ra
      -- 
    ra_3973_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1614_inst_ack_0, ack => convTransposeA_CP_3054_elements(111)); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	69 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (2) 
      -- CP-element group 112: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1611/phi_stmt_1611_sources/type_cast_1614/SplitProtocol/Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1611/phi_stmt_1611_sources/type_cast_1614/SplitProtocol/Update/ca
      -- 
    ca_3978_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1614_inst_ack_1, ack => convTransposeA_CP_3054_elements(112)); -- 
    -- CP-element group 113:  join  transition  output  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	111 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	120 
    -- CP-element group 113:  members (5) 
      -- CP-element group 113: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1611/$exit
      -- CP-element group 113: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1611/phi_stmt_1611_sources/$exit
      -- CP-element group 113: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1611/phi_stmt_1611_sources/type_cast_1614/$exit
      -- CP-element group 113: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1611/phi_stmt_1611_sources/type_cast_1614/SplitProtocol/$exit
      -- CP-element group 113: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1611/phi_stmt_1611_req
      -- 
    phi_stmt_1611_req_3979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1611_req_3979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(113), ack => phi_stmt_1611_req_0); -- 
    convTransposeA_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3054_elements(111) & convTransposeA_CP_3054_elements(112);
      gj_convTransposeA_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3054_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	69 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (2) 
      -- CP-element group 114: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/type_cast_1621/SplitProtocol/Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/type_cast_1621/SplitProtocol/Sample/ra
      -- 
    ra_3996_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1621_inst_ack_0, ack => convTransposeA_CP_3054_elements(114)); -- 
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	69 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/type_cast_1621/SplitProtocol/Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/type_cast_1621/SplitProtocol/Update/ca
      -- 
    ca_4001_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1621_inst_ack_1, ack => convTransposeA_CP_3054_elements(115)); -- 
    -- CP-element group 116:  join  transition  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	120 
    -- CP-element group 116:  members (5) 
      -- CP-element group 116: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1618/$exit
      -- CP-element group 116: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/$exit
      -- CP-element group 116: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/type_cast_1621/$exit
      -- CP-element group 116: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/type_cast_1621/SplitProtocol/$exit
      -- CP-element group 116: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1618/phi_stmt_1618_req
      -- 
    phi_stmt_1618_req_4002_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1618_req_4002_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(116), ack => phi_stmt_1618_req_0); -- 
    convTransposeA_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3054_elements(114) & convTransposeA_CP_3054_elements(115);
      gj_convTransposeA_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3054_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	69 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	119 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1627/SplitProtocol/Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1627/SplitProtocol/Sample/ra
      -- 
    ra_4019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1627_inst_ack_0, ack => convTransposeA_CP_3054_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	69 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (2) 
      -- CP-element group 118: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1627/SplitProtocol/Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1627/SplitProtocol/Update/ca
      -- 
    ca_4024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1627_inst_ack_1, ack => convTransposeA_CP_3054_elements(118)); -- 
    -- CP-element group 119:  join  transition  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	117 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (5) 
      -- CP-element group 119: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1624/$exit
      -- CP-element group 119: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/$exit
      -- CP-element group 119: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1627/$exit
      -- CP-element group 119: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1627/SplitProtocol/$exit
      -- CP-element group 119: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1624/phi_stmt_1624_req
      -- 
    phi_stmt_1624_req_4025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1624_req_4025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3054_elements(119), ack => phi_stmt_1624_req_0); -- 
    convTransposeA_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3054_elements(117) & convTransposeA_CP_3054_elements(118);
      gj_convTransposeA_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3054_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  join  transition  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	113 
    -- CP-element group 120: 	116 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_1293/ifx_xthen_ifx_xend123_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3054_elements(113) & convTransposeA_CP_3054_elements(116) & convTransposeA_CP_3054_elements(119);
      gj_convTransposeA_cp_element_group_120 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3054_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  merge  fork  transition  place  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	110 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121: 	123 
    -- CP-element group 121: 	124 
    -- CP-element group 121:  members (2) 
      -- CP-element group 121: 	 branch_block_stmt_1293/merge_stmt_1610_PhiReqMerge
      -- CP-element group 121: 	 branch_block_stmt_1293/merge_stmt_1610_PhiAck/$entry
      -- 
    convTransposeA_CP_3054_elements(121) <= OrReduce(convTransposeA_CP_3054_elements(110) & convTransposeA_CP_3054_elements(120));
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	125 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_1293/merge_stmt_1610_PhiAck/phi_stmt_1611_ack
      -- 
    phi_stmt_1611_ack_4030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1611_ack_0, ack => convTransposeA_CP_3054_elements(122)); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	121 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	125 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_1293/merge_stmt_1610_PhiAck/phi_stmt_1618_ack
      -- 
    phi_stmt_1618_ack_4031_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1618_ack_0, ack => convTransposeA_CP_3054_elements(123)); -- 
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	121 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	125 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_1293/merge_stmt_1610_PhiAck/phi_stmt_1624_ack
      -- 
    phi_stmt_1624_ack_4032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1624_ack_0, ack => convTransposeA_CP_3054_elements(124)); -- 
    -- CP-element group 125:  join  transition  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	122 
    -- CP-element group 125: 	123 
    -- CP-element group 125: 	124 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	1 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_1293/merge_stmt_1610_PhiAck/$exit
      -- 
    convTransposeA_cp_element_group_125: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_125"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3054_elements(122) & convTransposeA_CP_3054_elements(123) & convTransposeA_CP_3054_elements(124);
      gj_convTransposeA_cp_element_group_125 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3054_elements(125), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom81_1530_resized : std_logic_vector(13 downto 0);
    signal R_idxprom81_1530_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_1507_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_1507_scaled : std_logic_vector(13 downto 0);
    signal add41_1361 : std_logic_vector(15 downto 0);
    signal add54_1372 : std_logic_vector(15 downto 0);
    signal add73_1483 : std_logic_vector(63 downto 0);
    signal add75_1493 : std_logic_vector(63 downto 0);
    signal add86_1547 : std_logic_vector(31 downto 0);
    signal add93_1565 : std_logic_vector(15 downto 0);
    signal add_1345 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_1441 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1508_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1508_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1508_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1508_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1508_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1508_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1531_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1531_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1531_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1531_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1531_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1531_root_address : std_logic_vector(13 downto 0);
    signal arrayidx77_1510 : std_logic_vector(31 downto 0);
    signal arrayidx82_1533 : std_logic_vector(31 downto 0);
    signal call11_1314 : std_logic_vector(15 downto 0);
    signal call13_1317 : std_logic_vector(15 downto 0);
    signal call14_1320 : std_logic_vector(15 downto 0);
    signal call15_1323 : std_logic_vector(15 downto 0);
    signal call16_1336 : std_logic_vector(15 downto 0);
    signal call18_1348 : std_logic_vector(15 downto 0);
    signal call1_1299 : std_logic_vector(15 downto 0);
    signal call20_1351 : std_logic_vector(15 downto 0);
    signal call22_1354 : std_logic_vector(15 downto 0);
    signal call3_1302 : std_logic_vector(15 downto 0);
    signal call5_1305 : std_logic_vector(15 downto 0);
    signal call7_1308 : std_logic_vector(15 downto 0);
    signal call9_1311 : std_logic_vector(15 downto 0);
    signal call_1296 : std_logic_vector(15 downto 0);
    signal cmp101_1578 : std_logic_vector(0 downto 0);
    signal cmp112_1603 : std_logic_vector(0 downto 0);
    signal cmp_1552 : std_logic_vector(0 downto 0);
    signal conv107_1598 : std_logic_vector(31 downto 0);
    signal conv110_1393 : std_logic_vector(31 downto 0);
    signal conv17_1340 : std_logic_vector(31 downto 0);
    signal conv61_1465 : std_logic_vector(63 downto 0);
    signal conv64_1381 : std_logic_vector(63 downto 0);
    signal conv66_1469 : std_logic_vector(63 downto 0);
    signal conv69_1385 : std_logic_vector(63 downto 0);
    signal conv71_1473 : std_logic_vector(63 downto 0);
    signal conv85_1541 : std_logic_vector(31 downto 0);
    signal conv89_1389 : std_logic_vector(31 downto 0);
    signal conv_1327 : std_logic_vector(31 downto 0);
    signal idxprom81_1526 : std_logic_vector(63 downto 0);
    signal idxprom_1503 : std_logic_vector(63 downto 0);
    signal inc105_1582 : std_logic_vector(15 downto 0);
    signal inc105x_xinput_dim0x_x2_1587 : std_logic_vector(15 downto 0);
    signal inc_1573 : std_logic_vector(15 downto 0);
    signal indvar_1402 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_1636 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_1624 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_1423 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_1618 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_1416 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_1594 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_1611 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1409 : std_logic_vector(15 downto 0);
    signal mul50_1456 : std_logic_vector(15 downto 0);
    signal mul72_1478 : std_logic_vector(63 downto 0);
    signal mul74_1488 : std_logic_vector(63 downto 0);
    signal mul_1446 : std_logic_vector(15 downto 0);
    signal ptr_deref_1513_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1513_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1513_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1513_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1513_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1535_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1535_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1535_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1535_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1535_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1535_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_1333 : std_logic_vector(31 downto 0);
    signal shr111126_1399 : std_logic_vector(31 downto 0);
    signal shr80_1520 : std_logic_vector(63 downto 0);
    signal shr_1499 : std_logic_vector(31 downto 0);
    signal sub44_1451 : std_logic_vector(15 downto 0);
    signal sub57_1377 : std_logic_vector(15 downto 0);
    signal sub58_1461 : std_logic_vector(15 downto 0);
    signal sub_1366 : std_logic_vector(15 downto 0);
    signal tmp1_1436 : std_logic_vector(31 downto 0);
    signal tmp78_1514 : std_logic_vector(63 downto 0);
    signal type_cast_1331_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1359_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1370_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1397_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1406_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1408_wire : std_logic_vector(31 downto 0);
    signal type_cast_1413_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1415_wire : std_logic_vector(15 downto 0);
    signal type_cast_1420_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1422_wire : std_logic_vector(15 downto 0);
    signal type_cast_1427_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1429_wire : std_logic_vector(15 downto 0);
    signal type_cast_1434_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1497_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1518_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1524_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1545_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1563_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1571_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1591_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1614_wire : std_logic_vector(15 downto 0);
    signal type_cast_1617_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1621_wire : std_logic_vector(15 downto 0);
    signal type_cast_1623_wire : std_logic_vector(15 downto 0);
    signal type_cast_1627_wire : std_logic_vector(15 downto 0);
    signal type_cast_1629_wire : std_logic_vector(15 downto 0);
    signal type_cast_1634_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1642_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_1508_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1508_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1508_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1508_resized_base_address <= "00000000000000";
    array_obj_ref_1531_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1531_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1531_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1531_resized_base_address <= "00000000000000";
    ptr_deref_1513_word_offset_0 <= "00000000000000";
    ptr_deref_1535_word_offset_0 <= "00000000000000";
    type_cast_1331_wire_constant <= "00000000000000000000000000010000";
    type_cast_1359_wire_constant <= "1111111111111111";
    type_cast_1370_wire_constant <= "1111111111111111";
    type_cast_1397_wire_constant <= "00000000000000000000000000000010";
    type_cast_1406_wire_constant <= "00000000000000000000000000000000";
    type_cast_1413_wire_constant <= "0000000000000000";
    type_cast_1420_wire_constant <= "0000000000000000";
    type_cast_1427_wire_constant <= "0000000000000000";
    type_cast_1434_wire_constant <= "00000000000000000000000000000100";
    type_cast_1497_wire_constant <= "00000000000000000000000000000010";
    type_cast_1518_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1524_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_1545_wire_constant <= "00000000000000000000000000000100";
    type_cast_1563_wire_constant <= "0000000000000100";
    type_cast_1571_wire_constant <= "0000000000000001";
    type_cast_1591_wire_constant <= "0000000000000000";
    type_cast_1617_wire_constant <= "0000000000000000";
    type_cast_1634_wire_constant <= "00000000000000000000000000000001";
    type_cast_1642_wire_constant <= "0000000000000001";
    phi_stmt_1402: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1406_wire_constant & type_cast_1408_wire;
      req <= phi_stmt_1402_req_0 & phi_stmt_1402_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1402",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1402_ack_0,
          idata => idata,
          odata => indvar_1402,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1402
    phi_stmt_1409: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1413_wire_constant & type_cast_1415_wire;
      req <= phi_stmt_1409_req_0 & phi_stmt_1409_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1409",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1409_ack_0,
          idata => idata,
          odata => input_dim2x_x1_1409,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1409
    phi_stmt_1416: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1420_wire_constant & type_cast_1422_wire;
      req <= phi_stmt_1416_req_0 & phi_stmt_1416_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1416",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1416_ack_0,
          idata => idata,
          odata => input_dim1x_x1_1416,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1416
    phi_stmt_1423: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1427_wire_constant & type_cast_1429_wire;
      req <= phi_stmt_1423_req_0 & phi_stmt_1423_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1423",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1423_ack_0,
          idata => idata,
          odata => input_dim0x_x2_1423,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1423
    phi_stmt_1611: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1614_wire & type_cast_1617_wire_constant;
      req <= phi_stmt_1611_req_0 & phi_stmt_1611_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1611",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1611_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_1611,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1611
    phi_stmt_1618: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1621_wire & type_cast_1623_wire;
      req <= phi_stmt_1618_req_0 & phi_stmt_1618_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1618",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1618_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_1618,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1618
    phi_stmt_1624: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1627_wire & type_cast_1629_wire;
      req <= phi_stmt_1624_req_0 & phi_stmt_1624_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1624",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1624_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_1624,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1624
    -- flow-through select operator MUX_1593_inst
    input_dim1x_x2_1594 <= type_cast_1591_wire_constant when (cmp101_1578(0) /=  '0') else inc_1573;
    addr_of_1509_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1509_final_reg_req_0;
      addr_of_1509_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1509_final_reg_req_1;
      addr_of_1509_final_reg_ack_1<= rack(0);
      addr_of_1509_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1509_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1508_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx77_1510,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1532_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1532_final_reg_req_0;
      addr_of_1532_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1532_final_reg_req_1;
      addr_of_1532_final_reg_ack_1<= rack(0);
      addr_of_1532_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1532_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1531_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx82_1533,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1326_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1326_inst_req_0;
      type_cast_1326_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1326_inst_req_1;
      type_cast_1326_inst_ack_1<= rack(0);
      type_cast_1326_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1326_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_1323,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1327,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1339_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1339_inst_req_0;
      type_cast_1339_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1339_inst_req_1;
      type_cast_1339_inst_ack_1<= rack(0);
      type_cast_1339_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1339_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_1336,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_1340,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1380_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1380_inst_req_0;
      type_cast_1380_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1380_inst_req_1;
      type_cast_1380_inst_ack_1<= rack(0);
      type_cast_1380_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1380_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_1354,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv64_1381,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1384_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1384_inst_req_0;
      type_cast_1384_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1384_inst_req_1;
      type_cast_1384_inst_ack_1<= rack(0);
      type_cast_1384_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1384_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_1351,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv69_1385,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1388_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1388_inst_req_0;
      type_cast_1388_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1388_inst_req_1;
      type_cast_1388_inst_ack_1<= rack(0);
      type_cast_1388_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1388_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_1302,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv89_1389,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1392_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1392_inst_req_0;
      type_cast_1392_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1392_inst_req_1;
      type_cast_1392_inst_ack_1<= rack(0);
      type_cast_1392_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1392_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1296,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv110_1393,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1408_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1408_inst_req_0;
      type_cast_1408_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1408_inst_req_1;
      type_cast_1408_inst_ack_1<= rack(0);
      type_cast_1408_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1408_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1636,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1408_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1415_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1415_inst_req_0;
      type_cast_1415_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1415_inst_req_1;
      type_cast_1415_inst_ack_1<= rack(0);
      type_cast_1415_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1415_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_1611,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1415_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1422_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1422_inst_req_0;
      type_cast_1422_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1422_inst_req_1;
      type_cast_1422_inst_ack_1<= rack(0);
      type_cast_1422_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1422_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_1618,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1422_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1429_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1429_inst_req_0;
      type_cast_1429_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1429_inst_req_1;
      type_cast_1429_inst_ack_1<= rack(0);
      type_cast_1429_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1429_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_1624,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1429_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1464_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1464_inst_req_0;
      type_cast_1464_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1464_inst_req_1;
      type_cast_1464_inst_ack_1<= rack(0);
      type_cast_1464_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1464_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1409,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv61_1465,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1468_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1468_inst_req_0;
      type_cast_1468_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1468_inst_req_1;
      type_cast_1468_inst_ack_1<= rack(0);
      type_cast_1468_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1468_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub58_1461,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv66_1469,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1472_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1472_inst_req_0;
      type_cast_1472_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1472_inst_req_1;
      type_cast_1472_inst_ack_1<= rack(0);
      type_cast_1472_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1472_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub44_1451,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv71_1473,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1502_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1502_inst_req_0;
      type_cast_1502_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1502_inst_req_1;
      type_cast_1502_inst_ack_1<= rack(0);
      type_cast_1502_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1502_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr_1499,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_1503,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1540_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1540_inst_req_0;
      type_cast_1540_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1540_inst_req_1;
      type_cast_1540_inst_ack_1<= rack(0);
      type_cast_1540_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1540_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1409,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv85_1541,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1581_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1581_inst_req_0;
      type_cast_1581_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1581_inst_req_1;
      type_cast_1581_inst_ack_1<= rack(0);
      type_cast_1581_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1581_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp101_1578,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc105_1582,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1597_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1597_inst_req_0;
      type_cast_1597_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1597_inst_req_1;
      type_cast_1597_inst_ack_1<= rack(0);
      type_cast_1597_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1597_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc105x_xinput_dim0x_x2_1587,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv107_1598,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1614_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1614_inst_req_0;
      type_cast_1614_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1614_inst_req_1;
      type_cast_1614_inst_ack_1<= rack(0);
      type_cast_1614_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1614_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add93_1565,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1614_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1621_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1621_inst_req_0;
      type_cast_1621_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1621_inst_req_1;
      type_cast_1621_inst_ack_1<= rack(0);
      type_cast_1621_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1621_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_1416,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1621_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1623_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1623_inst_req_0;
      type_cast_1623_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1623_inst_req_1;
      type_cast_1623_inst_ack_1<= rack(0);
      type_cast_1623_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1623_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_1594,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1623_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1627_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1627_inst_req_0;
      type_cast_1627_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1627_inst_req_1;
      type_cast_1627_inst_ack_1<= rack(0);
      type_cast_1627_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1627_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_1423,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1627_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1629_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1629_inst_req_0;
      type_cast_1629_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1629_inst_req_1;
      type_cast_1629_inst_ack_1<= rack(0);
      type_cast_1629_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1629_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc105x_xinput_dim0x_x2_1587,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1629_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1508_index_1_rename
    process(R_idxprom_1507_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_1507_resized;
      ov(13 downto 0) := iv;
      R_idxprom_1507_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1508_index_1_resize
    process(idxprom_1503) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_1503;
      ov := iv(13 downto 0);
      R_idxprom_1507_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1508_root_address_inst
    process(array_obj_ref_1508_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1508_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1508_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1531_index_1_rename
    process(R_idxprom81_1530_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom81_1530_resized;
      ov(13 downto 0) := iv;
      R_idxprom81_1530_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1531_index_1_resize
    process(idxprom81_1526) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom81_1526;
      ov := iv(13 downto 0);
      R_idxprom81_1530_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1531_root_address_inst
    process(array_obj_ref_1531_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1531_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1531_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1513_addr_0
    process(ptr_deref_1513_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1513_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1513_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1513_base_resize
    process(arrayidx77_1510) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx77_1510;
      ov := iv(13 downto 0);
      ptr_deref_1513_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1513_gather_scatter
    process(ptr_deref_1513_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1513_data_0;
      ov(63 downto 0) := iv;
      tmp78_1514 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1513_root_address_inst
    process(ptr_deref_1513_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1513_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1513_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1535_addr_0
    process(ptr_deref_1535_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1535_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1535_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1535_base_resize
    process(arrayidx82_1533) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx82_1533;
      ov := iv(13 downto 0);
      ptr_deref_1535_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1535_gather_scatter
    process(tmp78_1514) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp78_1514;
      ov(63 downto 0) := iv;
      ptr_deref_1535_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1535_root_address_inst
    process(ptr_deref_1535_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1535_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1535_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1553_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_1552;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1553_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1553_branch_req_0,
          ack0 => if_stmt_1553_branch_ack_0,
          ack1 => if_stmt_1553_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1604_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp112_1603;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1604_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1604_branch_req_0,
          ack0 => if_stmt_1604_branch_ack_0,
          ack1 => if_stmt_1604_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1360_inst
    process(call7_1308) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_1308, type_cast_1359_wire_constant, tmp_var);
      add41_1361 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1371_inst
    process(call9_1311) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_1311, type_cast_1370_wire_constant, tmp_var);
      add54_1372 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1450_inst
    process(sub_1366, mul_1446) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_1366, mul_1446, tmp_var);
      sub44_1451 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1460_inst
    process(sub57_1377, mul50_1456) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub57_1377, mul50_1456, tmp_var);
      sub58_1461 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1564_inst
    process(input_dim2x_x1_1409) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_1409, type_cast_1563_wire_constant, tmp_var);
      add93_1565 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1572_inst
    process(input_dim1x_x1_1416) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_1416, type_cast_1571_wire_constant, tmp_var);
      inc_1573 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1586_inst
    process(inc105_1582, input_dim0x_x2_1423) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc105_1582, input_dim0x_x2_1423, tmp_var);
      inc105x_xinput_dim0x_x2_1587 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1440_inst
    process(add_1345, tmp1_1436) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_1345, tmp1_1436, tmp_var);
      add_src_0x_x0_1441 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1546_inst
    process(conv85_1541) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv85_1541, type_cast_1545_wire_constant, tmp_var);
      add86_1547 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1635_inst
    process(indvar_1402) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1402, type_cast_1634_wire_constant, tmp_var);
      indvarx_xnext_1636 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1482_inst
    process(mul72_1478, conv66_1469) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul72_1478, conv66_1469, tmp_var);
      add73_1483 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1492_inst
    process(mul74_1488, conv61_1465) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul74_1488, conv61_1465, tmp_var);
      add75_1493 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1525_inst
    process(shr80_1520) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr80_1520, type_cast_1524_wire_constant, tmp_var);
      idxprom81_1526 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1577_inst
    process(inc_1573, call1_1299) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_1573, call1_1299, tmp_var);
      cmp101_1578 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1602_inst
    process(conv107_1598, shr111126_1399) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv107_1598, shr111126_1399, tmp_var);
      cmp112_1603 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1398_inst
    process(conv110_1393) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv110_1393, type_cast_1397_wire_constant, tmp_var);
      shr111126_1399 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1498_inst
    process(add_src_0x_x0_1441) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_1441, type_cast_1497_wire_constant, tmp_var);
      shr_1499 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1519_inst
    process(add75_1493) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add75_1493, type_cast_1518_wire_constant, tmp_var);
      shr80_1520 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1445_inst
    process(input_dim0x_x2_1423, call13_1317) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x2_1423, call13_1317, tmp_var);
      mul_1446 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1455_inst
    process(input_dim1x_x1_1416, call13_1317) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_1416, call13_1317, tmp_var);
      mul50_1456 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1435_inst
    process(indvar_1402) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_1402, type_cast_1434_wire_constant, tmp_var);
      tmp1_1436 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1477_inst
    process(conv71_1473, conv69_1385) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv71_1473, conv69_1385, tmp_var);
      mul72_1478 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1487_inst
    process(add73_1483, conv64_1381) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add73_1483, conv64_1381, tmp_var);
      mul74_1488 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1344_inst
    process(shl_1333, conv17_1340) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_1333, conv17_1340, tmp_var);
      add_1345 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1332_inst
    process(conv_1327) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_1327, type_cast_1331_wire_constant, tmp_var);
      shl_1333 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1365_inst
    process(add41_1361, call14_1320) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add41_1361, call14_1320, tmp_var);
      sub_1366 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1376_inst
    process(add54_1372, call14_1320) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add54_1372, call14_1320, tmp_var);
      sub57_1377 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1551_inst
    process(add86_1547, conv89_1389) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add86_1547, conv89_1389, tmp_var);
      cmp_1552 <= tmp_var; --
    end process;
    -- shared split operator group (28) : array_obj_ref_1508_index_offset 
    ApIntAdd_group_28: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_1507_scaled;
      array_obj_ref_1508_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1508_index_offset_req_0;
      array_obj_ref_1508_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1508_index_offset_req_1;
      array_obj_ref_1508_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_28_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_28_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : array_obj_ref_1531_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom81_1530_scaled;
      array_obj_ref_1531_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1531_index_offset_req_0;
      array_obj_ref_1531_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1531_index_offset_req_1;
      array_obj_ref_1531_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared load operator group (0) : ptr_deref_1513_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1513_load_0_req_0;
      ptr_deref_1513_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1513_load_0_req_1;
      ptr_deref_1513_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1513_word_address_0;
      ptr_deref_1513_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_1535_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1535_store_0_req_0;
      ptr_deref_1535_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1535_store_0_req_1;
      ptr_deref_1535_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1535_word_address_0;
      data_in <= ptr_deref_1535_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block0_start_1347_inst RPIPE_Block0_start_1350_inst RPIPE_Block0_start_1353_inst RPIPE_Block0_start_1335_inst RPIPE_Block0_start_1322_inst RPIPE_Block0_start_1319_inst RPIPE_Block0_start_1316_inst RPIPE_Block0_start_1313_inst RPIPE_Block0_start_1310_inst RPIPE_Block0_start_1307_inst RPIPE_Block0_start_1304_inst RPIPE_Block0_start_1301_inst RPIPE_Block0_start_1298_inst RPIPE_Block0_start_1295_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block0_start_1347_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block0_start_1350_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block0_start_1353_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block0_start_1335_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block0_start_1322_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block0_start_1319_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block0_start_1316_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block0_start_1313_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block0_start_1310_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block0_start_1307_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block0_start_1304_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block0_start_1301_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block0_start_1298_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block0_start_1295_inst_req_0;
      RPIPE_Block0_start_1347_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block0_start_1350_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block0_start_1353_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block0_start_1335_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block0_start_1322_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block0_start_1319_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block0_start_1316_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block0_start_1313_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block0_start_1310_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block0_start_1307_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block0_start_1304_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block0_start_1301_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block0_start_1298_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block0_start_1295_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block0_start_1347_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block0_start_1350_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block0_start_1353_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block0_start_1335_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block0_start_1322_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block0_start_1319_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block0_start_1316_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block0_start_1313_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block0_start_1310_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block0_start_1307_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block0_start_1304_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block0_start_1301_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block0_start_1298_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block0_start_1295_inst_req_1;
      RPIPE_Block0_start_1347_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block0_start_1350_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block0_start_1353_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block0_start_1335_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block0_start_1322_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block0_start_1319_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block0_start_1316_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block0_start_1313_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block0_start_1310_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block0_start_1307_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block0_start_1304_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block0_start_1301_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block0_start_1298_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block0_start_1295_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call18_1348 <= data_out(223 downto 208);
      call20_1351 <= data_out(207 downto 192);
      call22_1354 <= data_out(191 downto 176);
      call16_1336 <= data_out(175 downto 160);
      call15_1323 <= data_out(159 downto 144);
      call14_1320 <= data_out(143 downto 128);
      call13_1317 <= data_out(127 downto 112);
      call11_1314 <= data_out(111 downto 96);
      call9_1311 <= data_out(95 downto 80);
      call7_1308 <= data_out(79 downto 64);
      call5_1305 <= data_out(63 downto 48);
      call3_1302 <= data_out(47 downto 32);
      call1_1299 <= data_out(31 downto 16);
      call_1296 <= data_out(15 downto 0);
      Block0_start_read_0_gI: SplitGuardInterface generic map(name => "Block0_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_start_read_0: InputPortRevised -- 
        generic map ( name => "Block0_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_start_pipe_read_req(0),
          oack => Block0_start_pipe_read_ack(0),
          odata => Block0_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block0_done_1640_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block0_done_1640_inst_req_0;
      WPIPE_Block0_done_1640_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block0_done_1640_inst_req_1;
      WPIPE_Block0_done_1640_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_1642_wire_constant;
      Block0_done_write_0_gI: SplitGuardInterface generic map(name => "Block0_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_done_pipe_write_req(0),
          oack => Block0_done_pipe_write_ack(0),
          odata => Block0_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeA_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    c : out  std_logic_vector(63 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal c_buffer :  std_logic_vector(63 downto 0);
  signal c_update_enable: Boolean;
  signal timer_CP_0_start: Boolean;
  signal timer_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal LOAD_count_22_load_0_req_0 : boolean;
  signal LOAD_count_22_load_0_ack_0 : boolean;
  signal LOAD_count_22_load_0_req_1 : boolean;
  signal LOAD_count_22_load_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= c_buffer;
  c <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_0: Block -- control-path 
    signal timer_CP_0_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    timer_CP_0_elements(0) <= timer_CP_0_start;
    timer_CP_0_symbol <= timer_CP_0_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_23/LOAD_count_22_sample_start_
      -- CP-element group 0: 	 assign_stmt_23/$entry
      -- CP-element group 0: 	 assign_stmt_23/LOAD_count_22_update_start_
      -- CP-element group 0: 	 assign_stmt_23/LOAD_count_22_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_23/LOAD_count_22_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_23/LOAD_count_22_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_23/LOAD_count_22_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_23/LOAD_count_22_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_23/LOAD_count_22_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_23/LOAD_count_22_Update/$entry
      -- CP-element group 0: 	 assign_stmt_23/LOAD_count_22_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_23/LOAD_count_22_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_23/LOAD_count_22_Update/word_access_complete/word_0/cr
      -- 
    cr_32_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_32_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => LOAD_count_22_load_0_req_1); -- 
    rr_21_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_21_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => LOAD_count_22_load_0_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 assign_stmt_23/LOAD_count_22_sample_completed_
      -- CP-element group 1: 	 assign_stmt_23/LOAD_count_22_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_23/LOAD_count_22_Sample/word_access_start/$exit
      -- CP-element group 1: 	 assign_stmt_23/LOAD_count_22_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 assign_stmt_23/LOAD_count_22_Sample/word_access_start/word_0/ra
      -- 
    ra_22_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_22_load_0_ack_0, ack => timer_CP_0_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_23/$exit
      -- CP-element group 2: 	 assign_stmt_23/LOAD_count_22_update_completed_
      -- CP-element group 2: 	 assign_stmt_23/LOAD_count_22_Update/$exit
      -- CP-element group 2: 	 assign_stmt_23/LOAD_count_22_Update/word_access_complete/$exit
      -- CP-element group 2: 	 assign_stmt_23/LOAD_count_22_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 assign_stmt_23/LOAD_count_22_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 assign_stmt_23/LOAD_count_22_Update/LOAD_count_22_Merge/$entry
      -- CP-element group 2: 	 assign_stmt_23/LOAD_count_22_Update/LOAD_count_22_Merge/$exit
      -- CP-element group 2: 	 assign_stmt_23/LOAD_count_22_Update/LOAD_count_22_Merge/merge_req
      -- CP-element group 2: 	 assign_stmt_23/LOAD_count_22_Update/LOAD_count_22_Merge/merge_ack
      -- 
    ca_33_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_22_load_0_ack_1, ack => timer_CP_0_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_count_22_data_0 : std_logic_vector(63 downto 0);
    signal LOAD_count_22_word_address_0 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    LOAD_count_22_word_address_0 <= "0";
    -- equivalence LOAD_count_22_gather_scatter
    process(LOAD_count_22_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_count_22_data_0;
      ov(63 downto 0) := iv;
      c_buffer <= ov(63 downto 0);
      --
    end process;
    -- shared load operator group (0) : LOAD_count_22_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_count_22_load_0_req_0;
      LOAD_count_22_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_count_22_load_0_req_1;
      LOAD_count_22_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_count_22_word_address_0;
      LOAD_count_22_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(0 downto 0),
          mtag => memory_space_0_lr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    ConvTranspose_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    ConvTranspose_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    ConvTranspose_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(17 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(10 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_3
  signal memory_space_3_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_3_lr_tag : std_logic_vector(17 downto 0);
  signal memory_space_3_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_3_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_3_sr_req :  std_logic_vector(1 downto 0);
  signal memory_space_3_sr_ack : std_logic_vector(1 downto 0);
  signal memory_space_3_sr_addr : std_logic_vector(27 downto 0);
  signal memory_space_3_sr_data : std_logic_vector(127 downto 0);
  signal memory_space_3_sr_tag : std_logic_vector(35 downto 0);
  signal memory_space_3_sc_req : std_logic_vector(1 downto 0);
  signal memory_space_3_sc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_3_sc_tag :  std_logic_vector(1 downto 0);
  -- declarations related to module convTranspose
  component convTranspose is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTranspose
  signal convTranspose_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTranspose_tag_out   : std_logic_vector(1 downto 0);
  signal convTranspose_start_req : std_logic;
  signal convTranspose_start_ack : std_logic;
  signal convTranspose_fin_req   : std_logic;
  signal convTranspose_fin_ack : std_logic;
  -- declarations related to module convTransposeA
  component convTransposeA is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeA
  signal convTransposeA_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeA_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeA_start_req : std_logic;
  signal convTransposeA_start_ack : std_logic;
  signal convTransposeA_fin_req   : std_logic;
  signal convTransposeA_fin_ack : std_logic;
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_c :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe Block0_done
  signal Block0_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_done
  signal Block0_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block0_start
  signal Block0_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_start
  signal Block0_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe ConvTranspose_input_pipe
  signal ConvTranspose_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe ConvTranspose_output_pipe
  signal ConvTranspose_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module convTranspose
  convTranspose_instance:convTranspose-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTranspose_start_req,
      start_ack => convTranspose_start_ack,
      fin_req => convTranspose_fin_req,
      fin_ack => convTranspose_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_3_lr_req => memory_space_3_lr_req(0 downto 0),
      memory_space_3_lr_ack => memory_space_3_lr_ack(0 downto 0),
      memory_space_3_lr_addr => memory_space_3_lr_addr(13 downto 0),
      memory_space_3_lr_tag => memory_space_3_lr_tag(17 downto 0),
      memory_space_3_lc_req => memory_space_3_lc_req(0 downto 0),
      memory_space_3_lc_ack => memory_space_3_lc_ack(0 downto 0),
      memory_space_3_lc_data => memory_space_3_lc_data(63 downto 0),
      memory_space_3_lc_tag => memory_space_3_lc_tag(0 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(17 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(0 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(10 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(63 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(0 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(0 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(1 downto 1),
      memory_space_3_sr_ack => memory_space_3_sr_ack(1 downto 1),
      memory_space_3_sr_addr => memory_space_3_sr_addr(27 downto 14),
      memory_space_3_sr_data => memory_space_3_sr_data(127 downto 64),
      memory_space_3_sr_tag => memory_space_3_sr_tag(35 downto 18),
      memory_space_3_sc_req => memory_space_3_sc_req(1 downto 1),
      memory_space_3_sc_ack => memory_space_3_sc_ack(1 downto 1),
      memory_space_3_sc_tag => memory_space_3_sc_tag(1 downto 1),
      Block0_done_pipe_read_req => Block0_done_pipe_read_req(0 downto 0),
      Block0_done_pipe_read_ack => Block0_done_pipe_read_ack(0 downto 0),
      Block0_done_pipe_read_data => Block0_done_pipe_read_data(15 downto 0),
      ConvTranspose_input_pipe_pipe_read_req => ConvTranspose_input_pipe_pipe_read_req(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_ack => ConvTranspose_input_pipe_pipe_read_ack(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_data => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
      ConvTranspose_output_pipe_pipe_write_req => ConvTranspose_output_pipe_pipe_write_req(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_ack => ConvTranspose_output_pipe_pipe_write_ack(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_data => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
      Block0_start_pipe_write_req => Block0_start_pipe_write_req(0 downto 0),
      Block0_start_pipe_write_ack => Block0_start_pipe_write_ack(0 downto 0),
      Block0_start_pipe_write_data => Block0_start_pipe_write_data(15 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      tag_in => convTranspose_tag_in,
      tag_out => convTranspose_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTranspose_tag_in <= (others => '0');
  convTranspose_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTranspose_start_req, start_ack => convTranspose_start_ack,  fin_req => convTranspose_fin_req,  fin_ack => convTranspose_fin_ack);
  -- module convTransposeA
  convTransposeA_instance:convTransposeA-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeA_start_req,
      start_ack => convTransposeA_start_ack,
      fin_req => convTransposeA_fin_req,
      fin_ack => convTransposeA_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(17 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(0 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(0 downto 0),
      memory_space_3_sr_ack => memory_space_3_sr_ack(0 downto 0),
      memory_space_3_sr_addr => memory_space_3_sr_addr(13 downto 0),
      memory_space_3_sr_data => memory_space_3_sr_data(63 downto 0),
      memory_space_3_sr_tag => memory_space_3_sr_tag(17 downto 0),
      memory_space_3_sc_req => memory_space_3_sc_req(0 downto 0),
      memory_space_3_sc_ack => memory_space_3_sc_ack(0 downto 0),
      memory_space_3_sc_tag => memory_space_3_sc_tag(0 downto 0),
      Block0_start_pipe_read_req => Block0_start_pipe_read_req(0 downto 0),
      Block0_start_pipe_read_ack => Block0_start_pipe_read_ack(0 downto 0),
      Block0_start_pipe_read_data => Block0_start_pipe_read_data(15 downto 0),
      Block0_done_pipe_write_req => Block0_done_pipe_write_req(0 downto 0),
      Block0_done_pipe_write_ack => Block0_done_pipe_write_ack(0 downto 0),
      Block0_done_pipe_write_data => Block0_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeA_tag_in,
      tag_out => convTransposeA_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeA_tag_in <= (others => '0');
  convTransposeA_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeA_start_req, start_ack => convTransposeA_start_ack,  fin_req => convTransposeA_fin_req,  fin_ack => convTransposeA_fin_ack);
  -- module timer
  timer_out_args <= timer_c ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      c => timer_c,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(0 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(0 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  Block0_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_done_pipe_read_req,
      read_ack => Block0_done_pipe_read_ack,
      read_data => Block0_done_pipe_read_data,
      write_req => Block0_done_pipe_write_req,
      write_ack => Block0_done_pipe_write_ack,
      write_data => Block0_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block0_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_start_pipe_read_req,
      read_ack => Block0_start_pipe_read_ack,
      read_data => Block0_start_pipe_read_data,
      write_req => Block0_start_pipe_write_req,
      write_ack => Block0_start_pipe_write_ack,
      write_data => Block0_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_input_pipe_pipe_read_req,
      read_ack => ConvTranspose_input_pipe_pipe_read_ack,
      read_data => ConvTranspose_input_pipe_pipe_read_data,
      write_req => ConvTranspose_input_pipe_pipe_write_req,
      write_ack => ConvTranspose_input_pipe_pipe_write_ack,
      write_data => ConvTranspose_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_output_pipe_pipe_read_req,
      read_ack => ConvTranspose_output_pipe_pipe_read_ack,
      read_data => ConvTranspose_output_pipe_pipe_read_data,
      write_req => ConvTranspose_output_pipe_pipe_write_req,
      write_ack => ConvTranspose_output_pipe_pipe_write_ack,
      write_data => ConvTranspose_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  dummyROM_memory_space_0: dummy_read_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      addr_width => 1,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_2: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_stores => 1,
      addr_width => 11,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_3: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_3",
      num_loads => 1,
      num_stores => 2,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_3_lr_addr,
      lr_req_in => memory_space_3_lr_req,
      lr_ack_out => memory_space_3_lr_ack,
      lr_tag_in => memory_space_3_lr_tag,
      lc_req_in => memory_space_3_lc_req,
      lc_ack_out => memory_space_3_lc_ack,
      lc_data_out => memory_space_3_lc_data,
      lc_tag_out => memory_space_3_lc_tag,
      sr_addr_in => memory_space_3_sr_addr,
      sr_data_in => memory_space_3_sr_data,
      sr_req_in => memory_space_3_sr_req,
      sr_ack_out => memory_space_3_sr_ack,
      sr_tag_in => memory_space_3_sr_tag,
      sc_req_in=> memory_space_3_sc_req,
      sc_ack_out => memory_space_3_sc_ack,
      sc_tag_out => memory_space_3_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
