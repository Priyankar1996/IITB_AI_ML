-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTranspose is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(10 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTranspose;
architecture convTranspose_arch of convTranspose is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTranspose_CP_39_start: Boolean;
  signal convTranspose_CP_39_symbol: Boolean;
  -- volatile/operator module components. 
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal type_cast_711_inst_req_0 : boolean;
  signal WPIPE_Block1_start_992_inst_req_0 : boolean;
  signal type_cast_711_inst_req_1 : boolean;
  signal type_cast_711_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_725_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1037_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_725_inst_ack_0 : boolean;
  signal type_cast_643_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_572_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_707_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1037_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1067_inst_ack_0 : boolean;
  signal type_cast_558_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_707_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1037_inst_ack_1 : boolean;
  signal type_cast_594_inst_req_0 : boolean;
  signal type_cast_711_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_725_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1037_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_725_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_48_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_48_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1028_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_572_inst_req_1 : boolean;
  signal type_cast_558_inst_req_1 : boolean;
  signal type_cast_643_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_572_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_518_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_518_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_572_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_518_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_518_inst_req_0 : boolean;
  signal type_cast_663_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_35_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_35_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_35_inst_req_1 : boolean;
  signal ptr_deref_602_store_0_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_35_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_689_inst_req_1 : boolean;
  signal WPIPE_Block0_start_983_inst_ack_1 : boolean;
  signal type_cast_643_inst_ack_1 : boolean;
  signal type_cast_39_inst_req_0 : boolean;
  signal type_cast_39_inst_ack_0 : boolean;
  signal type_cast_39_inst_req_1 : boolean;
  signal ptr_deref_602_store_0_req_0 : boolean;
  signal type_cast_39_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_135_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_135_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_554_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_135_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_135_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_554_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_48_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_48_inst_ack_1 : boolean;
  signal type_cast_52_inst_req_0 : boolean;
  signal type_cast_52_inst_ack_0 : boolean;
  signal type_cast_52_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1043_inst_req_1 : boolean;
  signal type_cast_52_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_60_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_60_inst_ack_0 : boolean;
  signal type_cast_558_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_60_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_60_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1058_inst_ack_1 : boolean;
  signal type_cast_643_inst_req_1 : boolean;
  signal type_cast_64_inst_req_0 : boolean;
  signal type_cast_64_inst_ack_0 : boolean;
  signal type_cast_64_inst_req_1 : boolean;
  signal type_cast_64_inst_ack_1 : boolean;
  signal addr_of_673_final_reg_ack_0 : boolean;
  signal type_cast_558_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_73_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_73_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1061_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_73_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_73_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1025_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1055_inst_ack_1 : boolean;
  signal type_cast_680_inst_ack_1 : boolean;
  signal type_cast_77_inst_req_0 : boolean;
  signal type_cast_77_inst_ack_0 : boolean;
  signal type_cast_77_inst_req_1 : boolean;
  signal type_cast_77_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_85_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_85_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_85_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1040_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_85_inst_ack_1 : boolean;
  signal type_cast_693_inst_ack_1 : boolean;
  signal type_cast_680_inst_req_1 : boolean;
  signal type_cast_89_inst_req_0 : boolean;
  signal type_cast_89_inst_ack_0 : boolean;
  signal type_cast_89_inst_req_1 : boolean;
  signal type_cast_89_inst_ack_1 : boolean;
  signal addr_of_673_final_reg_req_0 : boolean;
  signal if_stmt_1298_branch_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_98_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1040_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_98_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_98_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_98_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1046_inst_req_1 : boolean;
  signal type_cast_680_inst_ack_0 : boolean;
  signal type_cast_680_inst_req_0 : boolean;
  signal array_obj_ref_672_index_offset_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_689_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1016_inst_req_1 : boolean;
  signal type_cast_102_inst_req_0 : boolean;
  signal type_cast_102_inst_ack_0 : boolean;
  signal type_cast_102_inst_req_1 : boolean;
  signal type_cast_102_inst_ack_1 : boolean;
  signal addr_of_673_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_110_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_110_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_554_inst_ack_1 : boolean;
  signal addr_of_673_final_reg_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_110_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_110_inst_ack_1 : boolean;
  signal type_cast_693_inst_req_1 : boolean;
  signal array_obj_ref_672_index_offset_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_689_inst_req_0 : boolean;
  signal type_cast_114_inst_req_0 : boolean;
  signal type_cast_114_inst_ack_0 : boolean;
  signal type_cast_114_inst_req_1 : boolean;
  signal type_cast_114_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_992_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1025_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_554_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_123_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_123_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_123_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_123_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1067_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1016_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1046_inst_ack_1 : boolean;
  signal type_cast_127_inst_req_0 : boolean;
  signal type_cast_127_inst_ack_0 : boolean;
  signal type_cast_127_inst_req_1 : boolean;
  signal type_cast_127_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_707_inst_ack_1 : boolean;
  signal if_stmt_616_branch_ack_0 : boolean;
  signal WPIPE_Block1_start_992_inst_req_1 : boolean;
  signal type_cast_317_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1043_inst_req_0 : boolean;
  signal type_cast_317_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_986_inst_req_0 : boolean;
  signal type_cast_317_inst_req_1 : boolean;
  signal type_cast_317_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_326_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_326_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_995_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_326_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_326_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_995_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1281_inst_req_0 : boolean;
  signal type_cast_139_inst_req_0 : boolean;
  signal type_cast_139_inst_ack_0 : boolean;
  signal type_cast_139_inst_req_1 : boolean;
  signal type_cast_139_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1013_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_707_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_148_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1040_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_148_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_148_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_148_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1013_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1016_inst_req_0 : boolean;
  signal type_cast_152_inst_req_0 : boolean;
  signal type_cast_152_inst_ack_0 : boolean;
  signal type_cast_152_inst_req_1 : boolean;
  signal type_cast_152_inst_ack_1 : boolean;
  signal if_stmt_616_branch_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_160_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_160_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_160_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_160_inst_ack_1 : boolean;
  signal type_cast_693_inst_ack_0 : boolean;
  signal phi_stmt_453_ack_0 : boolean;
  signal type_cast_164_inst_req_0 : boolean;
  signal type_cast_164_inst_ack_0 : boolean;
  signal type_cast_164_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1040_inst_ack_1 : boolean;
  signal type_cast_164_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1061_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1013_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_590_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_173_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_173_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_173_inst_req_1 : boolean;
  signal WPIPE_Block0_start_980_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_173_inst_ack_1 : boolean;
  signal array_obj_ref_672_index_offset_ack_0 : boolean;
  signal WPIPE_Block1_start_1001_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_590_inst_req_1 : boolean;
  signal type_cast_177_inst_req_0 : boolean;
  signal type_cast_177_inst_ack_0 : boolean;
  signal type_cast_177_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1001_inst_ack_0 : boolean;
  signal type_cast_177_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_689_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_185_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_185_inst_ack_0 : boolean;
  signal type_cast_540_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_185_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_185_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_676_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_590_inst_ack_0 : boolean;
  signal type_cast_189_inst_req_0 : boolean;
  signal type_cast_189_inst_ack_0 : boolean;
  signal type_cast_189_inst_req_1 : boolean;
  signal type_cast_189_inst_ack_1 : boolean;
  signal type_cast_540_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_198_inst_req_0 : boolean;
  signal type_cast_910_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_198_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_198_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_198_inst_ack_1 : boolean;
  signal type_cast_693_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_676_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_590_inst_req_0 : boolean;
  signal type_cast_202_inst_req_0 : boolean;
  signal type_cast_202_inst_ack_0 : boolean;
  signal type_cast_202_inst_req_1 : boolean;
  signal type_cast_202_inst_ack_1 : boolean;
  signal type_cast_540_inst_ack_0 : boolean;
  signal type_cast_540_inst_req_0 : boolean;
  signal type_cast_211_inst_req_0 : boolean;
  signal type_cast_211_inst_ack_0 : boolean;
  signal type_cast_211_inst_req_1 : boolean;
  signal type_cast_211_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_980_inst_ack_0 : boolean;
  signal type_cast_215_inst_req_0 : boolean;
  signal type_cast_215_inst_ack_0 : boolean;
  signal type_cast_215_inst_req_1 : boolean;
  signal type_cast_215_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_980_inst_ack_1 : boolean;
  signal type_cast_219_inst_req_0 : boolean;
  signal type_cast_219_inst_ack_0 : boolean;
  signal type_cast_504_inst_ack_1 : boolean;
  signal type_cast_219_inst_req_1 : boolean;
  signal type_cast_219_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_536_inst_ack_1 : boolean;
  signal type_cast_233_inst_req_0 : boolean;
  signal type_cast_233_inst_ack_0 : boolean;
  signal type_cast_504_inst_req_1 : boolean;
  signal type_cast_233_inst_req_1 : boolean;
  signal type_cast_233_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_536_inst_req_1 : boolean;
  signal type_cast_237_inst_req_0 : boolean;
  signal type_cast_237_inst_ack_0 : boolean;
  signal type_cast_237_inst_req_1 : boolean;
  signal type_cast_237_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_536_inst_ack_0 : boolean;
  signal ptr_deref_602_store_0_ack_1 : boolean;
  signal type_cast_576_inst_ack_1 : boolean;
  signal type_cast_576_inst_req_1 : boolean;
  signal type_cast_241_inst_req_0 : boolean;
  signal type_cast_241_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1016_inst_ack_0 : boolean;
  signal type_cast_241_inst_req_1 : boolean;
  signal type_cast_241_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1028_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_536_inst_req_0 : boolean;
  signal ptr_deref_602_store_0_req_1 : boolean;
  signal type_cast_245_inst_req_0 : boolean;
  signal type_cast_245_inst_ack_0 : boolean;
  signal type_cast_504_inst_ack_0 : boolean;
  signal type_cast_245_inst_req_1 : boolean;
  signal type_cast_245_inst_ack_1 : boolean;
  signal if_stmt_616_branch_req_0 : boolean;
  signal WPIPE_Block1_start_992_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_263_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_263_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_263_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_263_inst_ack_1 : boolean;
  signal array_obj_ref_672_index_offset_req_0 : boolean;
  signal type_cast_576_inst_ack_0 : boolean;
  signal type_cast_576_inst_req_0 : boolean;
  signal type_cast_267_inst_req_0 : boolean;
  signal type_cast_267_inst_ack_0 : boolean;
  signal type_cast_267_inst_req_1 : boolean;
  signal type_cast_267_inst_ack_1 : boolean;
  signal type_cast_522_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_276_inst_req_0 : boolean;
  signal WPIPE_Block0_start_980_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_276_inst_ack_0 : boolean;
  signal type_cast_522_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_276_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_276_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_676_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_676_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1019_inst_req_0 : boolean;
  signal type_cast_280_inst_req_0 : boolean;
  signal type_cast_594_inst_ack_1 : boolean;
  signal type_cast_280_inst_ack_0 : boolean;
  signal type_cast_280_inst_req_1 : boolean;
  signal type_cast_280_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_288_inst_req_0 : boolean;
  signal type_cast_594_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_288_inst_ack_0 : boolean;
  signal type_cast_522_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_288_inst_req_1 : boolean;
  signal type_cast_910_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_288_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1019_inst_ack_0 : boolean;
  signal type_cast_292_inst_req_0 : boolean;
  signal type_cast_292_inst_ack_0 : boolean;
  signal type_cast_292_inst_req_1 : boolean;
  signal type_cast_292_inst_ack_1 : boolean;
  signal type_cast_522_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_301_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_301_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_301_inst_req_1 : boolean;
  signal type_cast_594_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_301_inst_ack_1 : boolean;
  signal type_cast_305_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1019_inst_req_1 : boolean;
  signal type_cast_305_inst_ack_0 : boolean;
  signal type_cast_305_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1019_inst_ack_1 : boolean;
  signal type_cast_305_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_313_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_313_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_313_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_313_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_995_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1052_inst_req_1 : boolean;
  signal WPIPE_Block1_start_995_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1052_inst_ack_1 : boolean;
  signal type_cast_330_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1281_inst_ack_0 : boolean;
  signal type_cast_330_inst_ack_0 : boolean;
  signal type_cast_330_inst_req_1 : boolean;
  signal type_cast_330_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_338_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1043_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_338_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_338_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_338_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_986_inst_ack_0 : boolean;
  signal type_cast_342_inst_req_0 : boolean;
  signal type_cast_342_inst_ack_0 : boolean;
  signal type_cast_342_inst_req_1 : boolean;
  signal type_cast_342_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1028_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1022_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_351_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_351_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_351_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_351_inst_ack_1 : boolean;
  signal type_cast_355_inst_req_0 : boolean;
  signal type_cast_355_inst_ack_0 : boolean;
  signal type_cast_355_inst_req_1 : boolean;
  signal type_cast_355_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1061_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_363_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_363_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_363_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_363_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1022_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_998_inst_req_0 : boolean;
  signal type_cast_367_inst_req_0 : boolean;
  signal type_cast_367_inst_ack_0 : boolean;
  signal type_cast_367_inst_req_1 : boolean;
  signal type_cast_367_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1001_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1061_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_998_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_376_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_376_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_376_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_376_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1064_inst_req_0 : boolean;
  signal type_cast_380_inst_req_0 : boolean;
  signal type_cast_380_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1001_inst_ack_1 : boolean;
  signal type_cast_380_inst_req_1 : boolean;
  signal type_cast_380_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1049_inst_req_0 : boolean;
  signal if_stmt_394_branch_req_0 : boolean;
  signal if_stmt_394_branch_ack_1 : boolean;
  signal if_stmt_394_branch_ack_0 : boolean;
  signal if_stmt_409_branch_req_0 : boolean;
  signal if_stmt_409_branch_ack_1 : boolean;
  signal if_stmt_409_branch_ack_0 : boolean;
  signal type_cast_436_inst_req_0 : boolean;
  signal type_cast_436_inst_ack_0 : boolean;
  signal type_cast_436_inst_req_1 : boolean;
  signal type_cast_436_inst_ack_1 : boolean;
  signal array_obj_ref_465_index_offset_req_0 : boolean;
  signal array_obj_ref_465_index_offset_ack_0 : boolean;
  signal array_obj_ref_465_index_offset_req_1 : boolean;
  signal array_obj_ref_465_index_offset_ack_1 : boolean;
  signal addr_of_466_final_reg_req_0 : boolean;
  signal addr_of_466_final_reg_ack_0 : boolean;
  signal addr_of_466_final_reg_req_1 : boolean;
  signal addr_of_466_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_469_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_469_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_469_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_469_inst_ack_1 : boolean;
  signal type_cast_473_inst_req_0 : boolean;
  signal type_cast_473_inst_ack_0 : boolean;
  signal type_cast_473_inst_req_1 : boolean;
  signal type_cast_473_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_482_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_482_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_482_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_482_inst_ack_1 : boolean;
  signal type_cast_486_inst_req_0 : boolean;
  signal type_cast_486_inst_ack_0 : boolean;
  signal type_cast_486_inst_req_1 : boolean;
  signal type_cast_486_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_500_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_500_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_500_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_500_inst_ack_1 : boolean;
  signal type_cast_504_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1013_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1058_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1055_inst_req_1 : boolean;
  signal type_cast_729_inst_req_0 : boolean;
  signal type_cast_729_inst_ack_0 : boolean;
  signal type_cast_729_inst_req_1 : boolean;
  signal type_cast_729_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1049_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_743_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_743_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_743_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_743_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1064_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1046_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1046_inst_req_0 : boolean;
  signal type_cast_747_inst_req_0 : boolean;
  signal type_cast_747_inst_ack_0 : boolean;
  signal type_cast_747_inst_req_1 : boolean;
  signal type_cast_747_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1049_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_761_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1034_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_761_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_761_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1034_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_761_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1064_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1058_inst_ack_0 : boolean;
  signal type_cast_765_inst_req_0 : boolean;
  signal type_cast_765_inst_ack_0 : boolean;
  signal type_cast_765_inst_req_1 : boolean;
  signal type_cast_765_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1067_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_989_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1010_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_779_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1034_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_779_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_989_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_779_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1034_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_779_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1058_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1010_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1055_inst_ack_0 : boolean;
  signal type_cast_783_inst_req_0 : boolean;
  signal type_cast_783_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1055_inst_req_0 : boolean;
  signal type_cast_783_inst_req_1 : boolean;
  signal type_cast_783_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1067_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1010_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_797_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_797_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1010_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_797_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_797_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_989_inst_ack_0 : boolean;
  signal type_cast_801_inst_req_0 : boolean;
  signal type_cast_801_inst_ack_0 : boolean;
  signal type_cast_801_inst_req_1 : boolean;
  signal type_cast_801_inst_ack_1 : boolean;
  signal phi_stmt_453_req_1 : boolean;
  signal WPIPE_Block2_start_1031_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1031_inst_req_1 : boolean;
  signal WPIPE_Block1_start_998_inst_ack_1 : boolean;
  signal ptr_deref_809_store_0_req_0 : boolean;
  signal ptr_deref_809_store_0_ack_0 : boolean;
  signal WPIPE_Block2_start_1025_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_983_inst_req_1 : boolean;
  signal WPIPE_Block1_start_998_inst_req_1 : boolean;
  signal ptr_deref_809_store_0_req_1 : boolean;
  signal WPIPE_Block1_start_1007_inst_ack_1 : boolean;
  signal ptr_deref_809_store_0_ack_1 : boolean;
  signal WPIPE_Block1_start_1007_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1052_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1052_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1025_inst_req_0 : boolean;
  signal if_stmt_823_branch_req_0 : boolean;
  signal WPIPE_Block1_start_1007_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_983_inst_ack_0 : boolean;
  signal if_stmt_823_branch_ack_1 : boolean;
  signal WPIPE_Block0_start_983_inst_req_0 : boolean;
  signal if_stmt_823_branch_ack_0 : boolean;
  signal WPIPE_Block2_start_1049_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1007_inst_req_0 : boolean;
  signal type_cast_834_inst_req_0 : boolean;
  signal type_cast_834_inst_ack_0 : boolean;
  signal type_cast_834_inst_req_1 : boolean;
  signal type_cast_834_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_989_inst_req_0 : boolean;
  signal type_cast_838_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1031_inst_ack_0 : boolean;
  signal type_cast_838_inst_ack_0 : boolean;
  signal type_cast_838_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1031_inst_req_0 : boolean;
  signal type_cast_838_inst_ack_1 : boolean;
  signal type_cast_842_inst_req_0 : boolean;
  signal type_cast_842_inst_ack_0 : boolean;
  signal type_cast_842_inst_req_1 : boolean;
  signal type_cast_842_inst_ack_1 : boolean;
  signal if_stmt_860_branch_req_0 : boolean;
  signal WPIPE_Block1_start_1004_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1022_inst_ack_1 : boolean;
  signal if_stmt_860_branch_ack_1 : boolean;
  signal if_stmt_860_branch_ack_0 : boolean;
  signal WPIPE_Block1_start_1022_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1004_inst_req_1 : boolean;
  signal type_cast_887_inst_req_0 : boolean;
  signal type_cast_887_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_977_inst_ack_1 : boolean;
  signal type_cast_887_inst_req_1 : boolean;
  signal type_cast_887_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_986_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1043_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_986_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1004_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1004_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1064_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_977_inst_req_1 : boolean;
  signal array_obj_ref_916_index_offset_req_0 : boolean;
  signal WPIPE_Block2_start_1028_inst_ack_1 : boolean;
  signal array_obj_ref_916_index_offset_ack_0 : boolean;
  signal array_obj_ref_916_index_offset_req_1 : boolean;
  signal array_obj_ref_916_index_offset_ack_1 : boolean;
  signal if_stmt_1298_branch_ack_0 : boolean;
  signal addr_of_917_final_reg_req_0 : boolean;
  signal addr_of_917_final_reg_ack_0 : boolean;
  signal addr_of_917_final_reg_req_1 : boolean;
  signal addr_of_917_final_reg_ack_1 : boolean;
  signal type_cast_1173_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1278_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1278_inst_ack_0 : boolean;
  signal type_cast_910_inst_req_1 : boolean;
  signal type_cast_910_inst_ack_1 : boolean;
  signal ptr_deref_920_store_0_req_0 : boolean;
  signal ptr_deref_920_store_0_ack_0 : boolean;
  signal ptr_deref_920_store_0_req_1 : boolean;
  signal ptr_deref_920_store_0_ack_1 : boolean;
  signal if_stmt_935_branch_req_0 : boolean;
  signal if_stmt_935_branch_ack_1 : boolean;
  signal type_cast_663_inst_req_0 : boolean;
  signal if_stmt_935_branch_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1281_inst_req_1 : boolean;
  signal call_stmt_946_call_req_0 : boolean;
  signal call_stmt_946_call_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1281_inst_ack_1 : boolean;
  signal call_stmt_946_call_req_1 : boolean;
  signal call_stmt_946_call_ack_1 : boolean;
  signal phi_stmt_1170_req_1 : boolean;
  signal type_cast_951_inst_req_0 : boolean;
  signal type_cast_951_inst_ack_0 : boolean;
  signal type_cast_663_inst_req_1 : boolean;
  signal type_cast_951_inst_req_1 : boolean;
  signal phi_stmt_660_req_1 : boolean;
  signal type_cast_951_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1278_inst_req_1 : boolean;
  signal phi_stmt_904_req_1 : boolean;
  signal WPIPE_Block0_start_953_inst_req_0 : boolean;
  signal WPIPE_Block0_start_953_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_953_inst_req_1 : boolean;
  signal WPIPE_Block0_start_953_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_956_inst_req_0 : boolean;
  signal WPIPE_Block0_start_956_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_956_inst_req_1 : boolean;
  signal WPIPE_Block0_start_956_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_959_inst_req_0 : boolean;
  signal WPIPE_Block0_start_959_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_959_inst_req_1 : boolean;
  signal WPIPE_Block0_start_959_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_962_inst_req_0 : boolean;
  signal WPIPE_Block0_start_962_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_962_inst_req_1 : boolean;
  signal WPIPE_Block0_start_962_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_965_inst_req_0 : boolean;
  signal WPIPE_Block0_start_965_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_965_inst_req_1 : boolean;
  signal WPIPE_Block0_start_965_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_968_inst_req_0 : boolean;
  signal WPIPE_Block0_start_968_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_968_inst_req_1 : boolean;
  signal WPIPE_Block0_start_968_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_971_inst_req_0 : boolean;
  signal WPIPE_Block0_start_971_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_971_inst_req_1 : boolean;
  signal WPIPE_Block0_start_971_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_974_inst_req_0 : boolean;
  signal WPIPE_Block0_start_974_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_974_inst_req_1 : boolean;
  signal WPIPE_Block0_start_974_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_977_inst_req_0 : boolean;
  signal WPIPE_Block0_start_977_inst_ack_0 : boolean;
  signal type_cast_459_inst_ack_1 : boolean;
  signal type_cast_459_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1070_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1070_inst_ack_0 : boolean;
  signal if_stmt_1298_branch_req_0 : boolean;
  signal WPIPE_Block3_start_1070_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1070_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1073_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1073_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1073_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1073_inst_ack_1 : boolean;
  signal type_cast_459_inst_ack_0 : boolean;
  signal type_cast_459_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1076_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1076_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1076_inst_req_1 : boolean;
  signal phi_stmt_904_req_0 : boolean;
  signal WPIPE_Block3_start_1076_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1079_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1079_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1079_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1079_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1082_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1082_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1082_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1082_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1085_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1085_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1085_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1085_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1088_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1088_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1284_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1088_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1088_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1091_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1091_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1284_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1091_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1091_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1094_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1094_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1094_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1094_inst_ack_1 : boolean;
  signal phi_stmt_453_req_0 : boolean;
  signal RPIPE_Block0_done_1098_inst_req_0 : boolean;
  signal RPIPE_Block0_done_1098_inst_ack_0 : boolean;
  signal RPIPE_Block0_done_1098_inst_req_1 : boolean;
  signal RPIPE_Block0_done_1098_inst_ack_1 : boolean;
  signal RPIPE_Block1_done_1101_inst_req_0 : boolean;
  signal RPIPE_Block1_done_1101_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1284_inst_ack_0 : boolean;
  signal RPIPE_Block1_done_1101_inst_req_1 : boolean;
  signal RPIPE_Block1_done_1101_inst_ack_1 : boolean;
  signal RPIPE_Block2_done_1104_inst_req_0 : boolean;
  signal RPIPE_Block2_done_1104_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1284_inst_req_0 : boolean;
  signal RPIPE_Block2_done_1104_inst_req_1 : boolean;
  signal RPIPE_Block2_done_1104_inst_ack_1 : boolean;
  signal RPIPE_Block3_done_1107_inst_req_0 : boolean;
  signal RPIPE_Block3_done_1107_inst_ack_0 : boolean;
  signal RPIPE_Block3_done_1107_inst_req_1 : boolean;
  signal RPIPE_Block3_done_1107_inst_ack_1 : boolean;
  signal call_stmt_1111_call_req_0 : boolean;
  signal call_stmt_1111_call_ack_0 : boolean;
  signal call_stmt_1111_call_req_1 : boolean;
  signal call_stmt_1111_call_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1275_inst_ack_1 : boolean;
  signal type_cast_1115_inst_req_0 : boolean;
  signal type_cast_1115_inst_ack_0 : boolean;
  signal type_cast_1115_inst_req_1 : boolean;
  signal type_cast_1115_inst_ack_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1122_inst_req_0 : boolean;
  signal WPIPE_elapsed_time_pipe_1122_inst_ack_0 : boolean;
  signal WPIPE_elapsed_time_pipe_1122_inst_req_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1122_inst_ack_1 : boolean;
  signal phi_stmt_1170_req_0 : boolean;
  signal if_stmt_1126_branch_req_0 : boolean;
  signal if_stmt_1126_branch_ack_1 : boolean;
  signal if_stmt_1126_branch_ack_0 : boolean;
  signal type_cast_1173_inst_ack_1 : boolean;
  signal type_cast_1153_inst_req_0 : boolean;
  signal type_cast_1153_inst_ack_0 : boolean;
  signal type_cast_1153_inst_req_1 : boolean;
  signal type_cast_1153_inst_ack_1 : boolean;
  signal type_cast_1173_inst_req_1 : boolean;
  signal phi_stmt_904_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1278_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1275_inst_req_1 : boolean;
  signal array_obj_ref_1182_index_offset_req_0 : boolean;
  signal array_obj_ref_1182_index_offset_ack_0 : boolean;
  signal array_obj_ref_1182_index_offset_req_1 : boolean;
  signal phi_stmt_660_ack_0 : boolean;
  signal array_obj_ref_1182_index_offset_ack_1 : boolean;
  signal type_cast_1173_inst_ack_0 : boolean;
  signal addr_of_1183_final_reg_req_0 : boolean;
  signal phi_stmt_660_req_0 : boolean;
  signal addr_of_1183_final_reg_ack_0 : boolean;
  signal phi_stmt_1170_ack_0 : boolean;
  signal addr_of_1183_final_reg_req_1 : boolean;
  signal type_cast_663_inst_ack_1 : boolean;
  signal addr_of_1183_final_reg_ack_1 : boolean;
  signal ptr_deref_1187_load_0_req_0 : boolean;
  signal ptr_deref_1187_load_0_ack_0 : boolean;
  signal ptr_deref_1187_load_0_req_1 : boolean;
  signal ptr_deref_1187_load_0_ack_1 : boolean;
  signal type_cast_1191_inst_req_0 : boolean;
  signal type_cast_1191_inst_ack_0 : boolean;
  signal type_cast_1191_inst_req_1 : boolean;
  signal type_cast_1191_inst_ack_1 : boolean;
  signal type_cast_1201_inst_req_0 : boolean;
  signal type_cast_1201_inst_ack_0 : boolean;
  signal type_cast_1201_inst_req_1 : boolean;
  signal type_cast_1201_inst_ack_1 : boolean;
  signal type_cast_1211_inst_req_0 : boolean;
  signal type_cast_1211_inst_ack_0 : boolean;
  signal type_cast_1211_inst_req_1 : boolean;
  signal type_cast_1211_inst_ack_1 : boolean;
  signal type_cast_1221_inst_req_0 : boolean;
  signal type_cast_1221_inst_ack_0 : boolean;
  signal type_cast_1221_inst_req_1 : boolean;
  signal type_cast_1221_inst_ack_1 : boolean;
  signal type_cast_1231_inst_req_0 : boolean;
  signal type_cast_1231_inst_ack_0 : boolean;
  signal type_cast_1231_inst_req_1 : boolean;
  signal type_cast_1231_inst_ack_1 : boolean;
  signal type_cast_1241_inst_req_0 : boolean;
  signal type_cast_1241_inst_ack_0 : boolean;
  signal type_cast_1241_inst_req_1 : boolean;
  signal type_cast_1241_inst_ack_1 : boolean;
  signal type_cast_1251_inst_req_0 : boolean;
  signal type_cast_1251_inst_ack_0 : boolean;
  signal type_cast_1251_inst_req_1 : boolean;
  signal type_cast_1251_inst_ack_1 : boolean;
  signal type_cast_1261_inst_req_0 : boolean;
  signal type_cast_1261_inst_ack_0 : boolean;
  signal type_cast_1261_inst_req_1 : boolean;
  signal type_cast_1261_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1263_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1263_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1263_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1263_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1266_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1266_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1266_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1266_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1269_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1269_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1269_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1269_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1272_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1272_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1272_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1272_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1275_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1275_inst_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTranspose_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTranspose_CP_39_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTranspose_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_39_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTranspose_CP_39_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_39_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTranspose_CP_39: Block -- control-path 
    signal convTranspose_CP_39_elements: BooleanArray(425 downto 0);
    -- 
  begin -- 
    convTranspose_CP_39_elements(0) <= convTranspose_CP_39_start;
    convTranspose_CP_39_symbol <= convTranspose_CP_39_elements(425);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	68 
    -- CP-element group 0: 	52 
    -- CP-element group 0: 	44 
    -- CP-element group 0: 	48 
    -- CP-element group 0: 	62 
    -- CP-element group 0: 	65 
    -- CP-element group 0: 	56 
    -- CP-element group 0: 	59 
    -- CP-element group 0: 	40 
    -- CP-element group 0: 	71 
    -- CP-element group 0: 	74 
    -- CP-element group 0: 	77 
    -- CP-element group 0: 	81 
    -- CP-element group 0: 	85 
    -- CP-element group 0: 	89 
    -- CP-element group 0: 	93 
    -- CP-element group 0: 	97 
    -- CP-element group 0: 	101 
    -- CP-element group 0: 	105 
    -- CP-element group 0: 	109 
    -- CP-element group 0: 	113 
    -- CP-element group 0: 	117 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	12 
    -- CP-element group 0: 	16 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	24 
    -- CP-element group 0: 	28 
    -- CP-element group 0: 	32 
    -- CP-element group 0: 	36 
    -- CP-element group 0:  members (101) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_33/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/branch_block_stmt_33__entry__
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393__entry__
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_35_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_35_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_35_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_39_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_39_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_39_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_139_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_52_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_52_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_52_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_64_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_64_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_64_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_77_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_77_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_77_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_89_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_89_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_89_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_102_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_102_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_102_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_114_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_114_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_114_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_127_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_127_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_127_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_317_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_317_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_139_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_139_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_152_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_152_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_152_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_164_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_305_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_164_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_164_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_177_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_177_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_177_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_189_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_189_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_189_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_202_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_202_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_202_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_211_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_211_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_211_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_215_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_215_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_215_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_219_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_219_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_219_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_233_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_233_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_233_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_237_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_237_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_237_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_241_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_241_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_241_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_245_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_245_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_245_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_267_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_267_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_267_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_280_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_280_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_280_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_292_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_292_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_292_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_305_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_305_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_317_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_330_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_330_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_330_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_342_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_342_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_342_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_355_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_355_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_355_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_367_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_367_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_367_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_380_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_380_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_380_Update/cr
      -- 
    rr_133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => RPIPE_ConvTranspose_input_pipe_35_inst_req_0); -- 
    cr_152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_39_inst_req_1); -- 
    cr_180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_52_inst_req_1); -- 
    cr_208_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_208_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_64_inst_req_1); -- 
    cr_236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_77_inst_req_1); -- 
    cr_264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_89_inst_req_1); -- 
    cr_292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_102_inst_req_1); -- 
    cr_320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_114_inst_req_1); -- 
    cr_348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_127_inst_req_1); -- 
    cr_754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_317_inst_req_1); -- 
    cr_376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_139_inst_req_1); -- 
    cr_404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_152_inst_req_1); -- 
    cr_432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_164_inst_req_1); -- 
    cr_460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_177_inst_req_1); -- 
    cr_488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_189_inst_req_1); -- 
    cr_516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_202_inst_req_1); -- 
    cr_530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_211_inst_req_1); -- 
    cr_544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_215_inst_req_1); -- 
    cr_558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_219_inst_req_1); -- 
    cr_572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_233_inst_req_1); -- 
    cr_586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_237_inst_req_1); -- 
    cr_600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_241_inst_req_1); -- 
    cr_614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_245_inst_req_1); -- 
    cr_642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_267_inst_req_1); -- 
    cr_670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_280_inst_req_1); -- 
    cr_698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_292_inst_req_1); -- 
    cr_726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_305_inst_req_1); -- 
    cr_782_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_782_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_330_inst_req_1); -- 
    cr_810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_342_inst_req_1); -- 
    cr_838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_355_inst_req_1); -- 
    cr_866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_367_inst_req_1); -- 
    cr_894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_380_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_35_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_35_update_start_
      -- CP-element group 1: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_35_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_35_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_35_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_35_Update/cr
      -- 
    ra_134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_35_inst_ack_0, ack => convTranspose_CP_39_elements(1)); -- 
    cr_138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(1), ack => RPIPE_ConvTranspose_input_pipe_35_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_48_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_48_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_48_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_35_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_35_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_35_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_39_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_39_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_39_Sample/rr
      -- 
    ca_139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_35_inst_ack_1, ack => convTranspose_CP_39_elements(2)); -- 
    rr_147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(2), ack => type_cast_39_inst_req_0); -- 
    rr_161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(2), ack => RPIPE_ConvTranspose_input_pipe_48_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_39_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_39_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_39_Sample/ra
      -- 
    ra_148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_39_inst_ack_0, ack => convTranspose_CP_39_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	57 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_39_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_39_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_39_Update/ca
      -- 
    ca_153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_39_inst_ack_1, ack => convTranspose_CP_39_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_48_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_48_update_start_
      -- CP-element group 5: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_48_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_48_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_48_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_48_Update/cr
      -- 
    ra_162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_48_inst_ack_0, ack => convTranspose_CP_39_elements(5)); -- 
    cr_166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(5), ack => RPIPE_ConvTranspose_input_pipe_48_inst_req_1); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_48_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_48_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_48_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_52_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_52_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_52_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_60_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_60_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_60_Sample/rr
      -- 
    ca_167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_48_inst_ack_1, ack => convTranspose_CP_39_elements(6)); -- 
    rr_175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(6), ack => type_cast_52_inst_req_0); -- 
    rr_189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(6), ack => RPIPE_ConvTranspose_input_pipe_60_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_52_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_52_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_52_Sample/ra
      -- 
    ra_176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_52_inst_ack_0, ack => convTranspose_CP_39_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	57 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_52_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_52_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_52_Update/ca
      -- 
    ca_181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_52_inst_ack_1, ack => convTranspose_CP_39_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_60_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_60_update_start_
      -- CP-element group 9: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_60_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_60_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_60_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_60_Update/cr
      -- 
    ra_190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_60_inst_ack_0, ack => convTranspose_CP_39_elements(9)); -- 
    cr_194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(9), ack => RPIPE_ConvTranspose_input_pipe_60_inst_req_1); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	13 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_60_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_60_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_60_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_64_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_64_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_64_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_73_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_73_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_73_Sample/rr
      -- 
    ca_195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_60_inst_ack_1, ack => convTranspose_CP_39_elements(10)); -- 
    rr_203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(10), ack => type_cast_64_inst_req_0); -- 
    rr_217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(10), ack => RPIPE_ConvTranspose_input_pipe_73_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_64_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_64_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_64_Sample/ra
      -- 
    ra_204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_64_inst_ack_0, ack => convTranspose_CP_39_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	60 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_64_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_64_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_64_Update/ca
      -- 
    ca_209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_64_inst_ack_1, ack => convTranspose_CP_39_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_73_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_73_update_start_
      -- CP-element group 13: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_73_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_73_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_73_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_73_Update/cr
      -- 
    ra_218_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_73_inst_ack_0, ack => convTranspose_CP_39_elements(13)); -- 
    cr_222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(13), ack => RPIPE_ConvTranspose_input_pipe_73_inst_req_1); -- 
    -- CP-element group 14:  fork  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_73_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_73_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_73_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_77_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_77_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_77_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_85_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_85_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_85_Sample/rr
      -- 
    ca_223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_73_inst_ack_1, ack => convTranspose_CP_39_elements(14)); -- 
    rr_231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(14), ack => type_cast_77_inst_req_0); -- 
    rr_245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(14), ack => RPIPE_ConvTranspose_input_pipe_85_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_77_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_77_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_77_Sample/ra
      -- 
    ra_232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_77_inst_ack_0, ack => convTranspose_CP_39_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	0 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	60 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_77_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_77_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_77_Update/ca
      -- 
    ca_237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_77_inst_ack_1, ack => convTranspose_CP_39_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_85_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_85_update_start_
      -- CP-element group 17: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_85_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_85_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_85_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_85_Update/cr
      -- 
    ra_246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_85_inst_ack_0, ack => convTranspose_CP_39_elements(17)); -- 
    cr_250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(17), ack => RPIPE_ConvTranspose_input_pipe_85_inst_req_1); -- 
    -- CP-element group 18:  fork  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18: 	21 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_85_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_85_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_85_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_89_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_89_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_89_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_98_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_98_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_98_Sample/rr
      -- 
    ca_251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_85_inst_ack_1, ack => convTranspose_CP_39_elements(18)); -- 
    rr_259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(18), ack => type_cast_89_inst_req_0); -- 
    rr_273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(18), ack => RPIPE_ConvTranspose_input_pipe_98_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_89_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_89_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_89_Sample/ra
      -- 
    ra_260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_89_inst_ack_0, ack => convTranspose_CP_39_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	63 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_89_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_89_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_89_Update/ca
      -- 
    ca_265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_89_inst_ack_1, ack => convTranspose_CP_39_elements(20)); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_98_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_98_update_start_
      -- CP-element group 21: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_98_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_98_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_98_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_98_Update/cr
      -- 
    ra_274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_98_inst_ack_0, ack => convTranspose_CP_39_elements(21)); -- 
    cr_278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(21), ack => RPIPE_ConvTranspose_input_pipe_98_inst_req_1); -- 
    -- CP-element group 22:  fork  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22: 	25 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_98_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_98_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_98_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_102_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_102_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_102_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_110_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_110_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_110_Sample/rr
      -- 
    ca_279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_98_inst_ack_1, ack => convTranspose_CP_39_elements(22)); -- 
    rr_287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(22), ack => type_cast_102_inst_req_0); -- 
    rr_301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(22), ack => RPIPE_ConvTranspose_input_pipe_110_inst_req_0); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_102_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_102_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_102_Sample/ra
      -- 
    ra_288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_102_inst_ack_0, ack => convTranspose_CP_39_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	0 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	63 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_102_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_102_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_102_Update/ca
      -- 
    ca_293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_102_inst_ack_1, ack => convTranspose_CP_39_elements(24)); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	22 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_110_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_110_update_start_
      -- CP-element group 25: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_110_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_110_Sample/ra
      -- CP-element group 25: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_110_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_110_Update/cr
      -- 
    ra_302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_110_inst_ack_0, ack => convTranspose_CP_39_elements(25)); -- 
    cr_306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(25), ack => RPIPE_ConvTranspose_input_pipe_110_inst_req_1); -- 
    -- CP-element group 26:  fork  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: 	29 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_110_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_110_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_110_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_114_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_114_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_114_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_123_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_123_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_123_Sample/rr
      -- 
    ca_307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_110_inst_ack_1, ack => convTranspose_CP_39_elements(26)); -- 
    rr_315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(26), ack => type_cast_114_inst_req_0); -- 
    rr_329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(26), ack => RPIPE_ConvTranspose_input_pipe_123_inst_req_0); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_114_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_114_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_114_Sample/ra
      -- 
    ra_316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_114_inst_ack_0, ack => convTranspose_CP_39_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	0 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	66 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_114_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_114_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_114_Update/ca
      -- 
    ca_321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_114_inst_ack_1, ack => convTranspose_CP_39_elements(28)); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	26 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_123_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_123_update_start_
      -- CP-element group 29: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_123_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_123_Sample/ra
      -- CP-element group 29: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_123_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_123_Update/cr
      -- 
    ra_330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_123_inst_ack_0, ack => convTranspose_CP_39_elements(29)); -- 
    cr_334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(29), ack => RPIPE_ConvTranspose_input_pipe_123_inst_req_1); -- 
    -- CP-element group 30:  fork  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: 	33 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_135_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_123_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_123_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_123_Update/ca
      -- CP-element group 30: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_127_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_127_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_127_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_135_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_135_Sample/$entry
      -- 
    ca_335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_123_inst_ack_1, ack => convTranspose_CP_39_elements(30)); -- 
    rr_343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(30), ack => type_cast_127_inst_req_0); -- 
    rr_357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(30), ack => RPIPE_ConvTranspose_input_pipe_135_inst_req_0); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_127_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_127_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_127_Sample/ra
      -- 
    ra_344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_127_inst_ack_0, ack => convTranspose_CP_39_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	0 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	66 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_127_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_127_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_127_Update/ca
      -- 
    ca_349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_127_inst_ack_1, ack => convTranspose_CP_39_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	30 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_135_Sample/ra
      -- CP-element group 33: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_135_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_135_Update/cr
      -- CP-element group 33: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_135_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_135_update_start_
      -- CP-element group 33: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_135_Sample/$exit
      -- 
    ra_358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_135_inst_ack_0, ack => convTranspose_CP_39_elements(33)); -- 
    cr_362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(33), ack => RPIPE_ConvTranspose_input_pipe_135_inst_req_1); -- 
    -- CP-element group 34:  fork  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	37 
    -- CP-element group 34:  members (9) 
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_135_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_135_Update/ca
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_139_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_135_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_139_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_139_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_148_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_148_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_148_Sample/rr
      -- 
    ca_363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_135_inst_ack_1, ack => convTranspose_CP_39_elements(34)); -- 
    rr_371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(34), ack => type_cast_139_inst_req_0); -- 
    rr_385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(34), ack => RPIPE_ConvTranspose_input_pipe_148_inst_req_0); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_139_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_139_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_139_Sample/ra
      -- 
    ra_372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_139_inst_ack_0, ack => convTranspose_CP_39_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	0 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	69 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_139_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_139_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_139_Update/ca
      -- 
    ca_377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_139_inst_ack_1, ack => convTranspose_CP_39_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_148_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_148_update_start_
      -- CP-element group 37: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_148_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_148_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_148_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_148_Update/cr
      -- 
    ra_386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_148_inst_ack_0, ack => convTranspose_CP_39_elements(37)); -- 
    cr_390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(37), ack => RPIPE_ConvTranspose_input_pipe_148_inst_req_1); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	41 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_148_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_148_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_148_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_152_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_152_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_152_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_160_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_160_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_160_Sample/rr
      -- 
    ca_391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_148_inst_ack_1, ack => convTranspose_CP_39_elements(38)); -- 
    rr_399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(38), ack => type_cast_152_inst_req_0); -- 
    rr_413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(38), ack => RPIPE_ConvTranspose_input_pipe_160_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_152_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_152_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_152_Sample/ra
      -- 
    ra_400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_152_inst_ack_0, ack => convTranspose_CP_39_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	0 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	69 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_152_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_152_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_152_Update/ca
      -- 
    ca_405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_152_inst_ack_1, ack => convTranspose_CP_39_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	38 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_160_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_160_update_start_
      -- CP-element group 41: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_160_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_160_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_160_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_160_Update/cr
      -- 
    ra_414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_160_inst_ack_0, ack => convTranspose_CP_39_elements(41)); -- 
    cr_418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(41), ack => RPIPE_ConvTranspose_input_pipe_160_inst_req_1); -- 
    -- CP-element group 42:  fork  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42: 	45 
    -- CP-element group 42:  members (9) 
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_160_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_160_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_160_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_164_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_164_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_164_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_173_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_173_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_173_Sample/rr
      -- 
    ca_419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_160_inst_ack_1, ack => convTranspose_CP_39_elements(42)); -- 
    rr_427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(42), ack => type_cast_164_inst_req_0); -- 
    rr_441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(42), ack => RPIPE_ConvTranspose_input_pipe_173_inst_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_164_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_164_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_164_Sample/ra
      -- 
    ra_428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_164_inst_ack_0, ack => convTranspose_CP_39_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	0 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	72 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_164_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_164_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_164_Update/ca
      -- 
    ca_433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_164_inst_ack_1, ack => convTranspose_CP_39_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	42 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_173_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_173_update_start_
      -- CP-element group 45: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_173_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_173_Sample/ra
      -- CP-element group 45: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_173_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_173_Update/cr
      -- 
    ra_442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_173_inst_ack_0, ack => convTranspose_CP_39_elements(45)); -- 
    cr_446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(45), ack => RPIPE_ConvTranspose_input_pipe_173_inst_req_1); -- 
    -- CP-element group 46:  fork  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46: 	49 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_173_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_173_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_173_Update/ca
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_177_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_177_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_177_Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_185_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_185_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_185_Sample/rr
      -- 
    ca_447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_173_inst_ack_1, ack => convTranspose_CP_39_elements(46)); -- 
    rr_469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(46), ack => RPIPE_ConvTranspose_input_pipe_185_inst_req_0); -- 
    rr_455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(46), ack => type_cast_177_inst_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_177_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_177_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_177_Sample/ra
      -- 
    ra_456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_177_inst_ack_0, ack => convTranspose_CP_39_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	0 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	72 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_177_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_177_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_177_Update/ca
      -- 
    ca_461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_177_inst_ack_1, ack => convTranspose_CP_39_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	46 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_185_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_185_update_start_
      -- CP-element group 49: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_185_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_185_Sample/ra
      -- CP-element group 49: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_185_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_185_Update/cr
      -- 
    ra_470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_185_inst_ack_0, ack => convTranspose_CP_39_elements(49)); -- 
    cr_474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(49), ack => RPIPE_ConvTranspose_input_pipe_185_inst_req_1); -- 
    -- CP-element group 50:  fork  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	53 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_185_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_185_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_185_Update/ca
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_189_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_189_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_189_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_198_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_198_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_198_Sample/rr
      -- 
    ca_475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_185_inst_ack_1, ack => convTranspose_CP_39_elements(50)); -- 
    rr_483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(50), ack => type_cast_189_inst_req_0); -- 
    rr_497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(50), ack => RPIPE_ConvTranspose_input_pipe_198_inst_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_189_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_189_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_189_Sample/ra
      -- 
    ra_484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_189_inst_ack_0, ack => convTranspose_CP_39_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	0 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	75 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_189_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_189_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_189_Update/ca
      -- 
    ca_489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_189_inst_ack_1, ack => convTranspose_CP_39_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	50 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (6) 
      -- CP-element group 53: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_198_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_198_update_start_
      -- CP-element group 53: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_198_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_198_Sample/ra
      -- CP-element group 53: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_198_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_198_Update/cr
      -- 
    ra_498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_198_inst_ack_0, ack => convTranspose_CP_39_elements(53)); -- 
    cr_502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(53), ack => RPIPE_ConvTranspose_input_pipe_198_inst_req_1); -- 
    -- CP-element group 54:  fork  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54: 	78 
    -- CP-element group 54:  members (9) 
      -- CP-element group 54: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_198_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_198_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_198_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_202_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_202_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_202_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_263_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_263_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_263_Sample/rr
      -- 
    ca_503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_198_inst_ack_1, ack => convTranspose_CP_39_elements(54)); -- 
    rr_511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(54), ack => type_cast_202_inst_req_0); -- 
    rr_623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(54), ack => RPIPE_ConvTranspose_input_pipe_263_inst_req_0); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_202_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_202_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_202_Sample/ra
      -- 
    ra_512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_202_inst_ack_0, ack => convTranspose_CP_39_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	0 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	75 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_202_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_202_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_202_Update/ca
      -- 
    ca_517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_202_inst_ack_1, ack => convTranspose_CP_39_elements(56)); -- 
    -- CP-element group 57:  join  transition  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	4 
    -- CP-element group 57: 	8 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_211_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_211_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_211_Sample/rr
      -- 
    rr_525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(57), ack => type_cast_211_inst_req_0); -- 
    convTranspose_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(4) & convTranspose_CP_39_elements(8);
      gj_convTranspose_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_211_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_211_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_211_Sample/ra
      -- 
    ra_526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_211_inst_ack_0, ack => convTranspose_CP_39_elements(58)); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	0 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	118 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_211_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_211_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_211_Update/ca
      -- 
    ca_531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_211_inst_ack_1, ack => convTranspose_CP_39_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	12 
    -- CP-element group 60: 	16 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_215_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_215_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_215_Sample/rr
      -- 
    rr_539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(60), ack => type_cast_215_inst_req_0); -- 
    convTranspose_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(12) & convTranspose_CP_39_elements(16);
      gj_convTranspose_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_215_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_215_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_215_Sample/ra
      -- 
    ra_540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_215_inst_ack_0, ack => convTranspose_CP_39_elements(61)); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	0 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	118 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_215_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_215_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_215_Update/ca
      -- 
    ca_545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_215_inst_ack_1, ack => convTranspose_CP_39_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	20 
    -- CP-element group 63: 	24 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_219_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_219_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_219_Sample/rr
      -- 
    rr_553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(63), ack => type_cast_219_inst_req_0); -- 
    convTranspose_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(20) & convTranspose_CP_39_elements(24);
      gj_convTranspose_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_219_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_219_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_219_Sample/ra
      -- 
    ra_554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_219_inst_ack_0, ack => convTranspose_CP_39_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	0 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	118 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_219_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_219_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_219_Update/ca
      -- 
    ca_559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_219_inst_ack_1, ack => convTranspose_CP_39_elements(65)); -- 
    -- CP-element group 66:  join  transition  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	28 
    -- CP-element group 66: 	32 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_233_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_233_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_233_Sample/rr
      -- 
    rr_567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(66), ack => type_cast_233_inst_req_0); -- 
    convTranspose_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(28) & convTranspose_CP_39_elements(32);
      gj_convTranspose_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_233_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_233_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_233_Sample/ra
      -- 
    ra_568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_233_inst_ack_0, ack => convTranspose_CP_39_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	0 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	118 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_233_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_233_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_233_Update/ca
      -- 
    ca_573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_233_inst_ack_1, ack => convTranspose_CP_39_elements(68)); -- 
    -- CP-element group 69:  join  transition  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	40 
    -- CP-element group 69: 	36 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_237_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_237_Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_237_Sample/rr
      -- 
    rr_581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(69), ack => type_cast_237_inst_req_0); -- 
    convTranspose_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(40) & convTranspose_CP_39_elements(36);
      gj_convTranspose_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_237_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_237_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_237_Sample/ra
      -- 
    ra_582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_237_inst_ack_0, ack => convTranspose_CP_39_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	0 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	118 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_237_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_237_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_237_Update/ca
      -- 
    ca_587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_237_inst_ack_1, ack => convTranspose_CP_39_elements(71)); -- 
    -- CP-element group 72:  join  transition  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	44 
    -- CP-element group 72: 	48 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_241_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_241_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_241_Sample/rr
      -- 
    rr_595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(72), ack => type_cast_241_inst_req_0); -- 
    convTranspose_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(44) & convTranspose_CP_39_elements(48);
      gj_convTranspose_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_241_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_241_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_241_Sample/ra
      -- 
    ra_596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_241_inst_ack_0, ack => convTranspose_CP_39_elements(73)); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	0 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	118 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_241_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_241_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_241_Update/ca
      -- 
    ca_601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_241_inst_ack_1, ack => convTranspose_CP_39_elements(74)); -- 
    -- CP-element group 75:  join  transition  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	52 
    -- CP-element group 75: 	56 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_245_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_245_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_245_Sample/rr
      -- 
    rr_609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(75), ack => type_cast_245_inst_req_0); -- 
    convTranspose_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(52) & convTranspose_CP_39_elements(56);
      gj_convTranspose_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_245_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_245_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_245_Sample/ra
      -- 
    ra_610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_245_inst_ack_0, ack => convTranspose_CP_39_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	0 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	118 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_245_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_245_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_245_Update/ca
      -- 
    ca_615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_245_inst_ack_1, ack => convTranspose_CP_39_elements(77)); -- 
    -- CP-element group 78:  transition  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	54 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (6) 
      -- CP-element group 78: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_263_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_263_update_start_
      -- CP-element group 78: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_263_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_263_Sample/ra
      -- CP-element group 78: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_263_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_263_Update/cr
      -- 
    ra_624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_263_inst_ack_0, ack => convTranspose_CP_39_elements(78)); -- 
    cr_628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(78), ack => RPIPE_ConvTranspose_input_pipe_263_inst_req_1); -- 
    -- CP-element group 79:  fork  transition  input  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79: 	82 
    -- CP-element group 79:  members (9) 
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_263_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_263_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_263_Update/ca
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_267_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_267_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_267_Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_276_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_276_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_276_Sample/rr
      -- 
    ca_629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_263_inst_ack_1, ack => convTranspose_CP_39_elements(79)); -- 
    rr_637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(79), ack => type_cast_267_inst_req_0); -- 
    rr_651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(79), ack => RPIPE_ConvTranspose_input_pipe_276_inst_req_0); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_267_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_267_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_267_Sample/ra
      -- 
    ra_638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_267_inst_ack_0, ack => convTranspose_CP_39_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	0 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	118 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_267_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_267_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_267_Update/ca
      -- 
    ca_643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_267_inst_ack_1, ack => convTranspose_CP_39_elements(81)); -- 
    -- CP-element group 82:  transition  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	79 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (6) 
      -- CP-element group 82: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_276_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_276_update_start_
      -- CP-element group 82: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_276_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_276_Sample/ra
      -- CP-element group 82: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_276_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_276_Update/cr
      -- 
    ra_652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_276_inst_ack_0, ack => convTranspose_CP_39_elements(82)); -- 
    cr_656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(82), ack => RPIPE_ConvTranspose_input_pipe_276_inst_req_1); -- 
    -- CP-element group 83:  fork  transition  input  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83: 	86 
    -- CP-element group 83:  members (9) 
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_276_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_276_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_276_Update/ca
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_280_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_280_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_280_Sample/rr
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_288_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_288_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_288_Sample/rr
      -- 
    ca_657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_276_inst_ack_1, ack => convTranspose_CP_39_elements(83)); -- 
    rr_665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(83), ack => type_cast_280_inst_req_0); -- 
    rr_679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(83), ack => RPIPE_ConvTranspose_input_pipe_288_inst_req_0); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_280_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_280_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_280_Sample/ra
      -- 
    ra_666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_280_inst_ack_0, ack => convTranspose_CP_39_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	0 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	118 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_280_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_280_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_280_Update/ca
      -- 
    ca_671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_280_inst_ack_1, ack => convTranspose_CP_39_elements(85)); -- 
    -- CP-element group 86:  transition  input  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	83 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (6) 
      -- CP-element group 86: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_288_sample_completed_
      -- CP-element group 86: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_288_update_start_
      -- CP-element group 86: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_288_Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_288_Sample/ra
      -- CP-element group 86: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_288_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_288_Update/cr
      -- 
    ra_680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_288_inst_ack_0, ack => convTranspose_CP_39_elements(86)); -- 
    cr_684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(86), ack => RPIPE_ConvTranspose_input_pipe_288_inst_req_1); -- 
    -- CP-element group 87:  fork  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87: 	90 
    -- CP-element group 87:  members (9) 
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_288_update_completed_
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_288_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_288_Update/ca
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_292_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_292_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_292_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_301_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_301_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_301_Sample/rr
      -- 
    ca_685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_288_inst_ack_1, ack => convTranspose_CP_39_elements(87)); -- 
    rr_693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(87), ack => type_cast_292_inst_req_0); -- 
    rr_707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(87), ack => RPIPE_ConvTranspose_input_pipe_301_inst_req_0); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_292_sample_completed_
      -- CP-element group 88: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_292_Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_292_Sample/ra
      -- 
    ra_694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_292_inst_ack_0, ack => convTranspose_CP_39_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	0 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	118 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_292_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_292_Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_292_Update/ca
      -- 
    ca_699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_292_inst_ack_1, ack => convTranspose_CP_39_elements(89)); -- 
    -- CP-element group 90:  transition  input  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	87 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (6) 
      -- CP-element group 90: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_301_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_301_update_start_
      -- CP-element group 90: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_301_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_301_Sample/ra
      -- CP-element group 90: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_301_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_301_Update/cr
      -- 
    ra_708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_301_inst_ack_0, ack => convTranspose_CP_39_elements(90)); -- 
    cr_712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(90), ack => RPIPE_ConvTranspose_input_pipe_301_inst_req_1); -- 
    -- CP-element group 91:  fork  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91: 	94 
    -- CP-element group 91:  members (9) 
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_301_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_301_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_301_Update/ca
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_305_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_305_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_305_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_313_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_313_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_313_Sample/rr
      -- 
    ca_713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_301_inst_ack_1, ack => convTranspose_CP_39_elements(91)); -- 
    rr_721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(91), ack => type_cast_305_inst_req_0); -- 
    rr_735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(91), ack => RPIPE_ConvTranspose_input_pipe_313_inst_req_0); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_305_sample_completed_
      -- CP-element group 92: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_305_Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_305_Sample/ra
      -- 
    ra_722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_305_inst_ack_0, ack => convTranspose_CP_39_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	0 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	118 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_305_Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_305_update_completed_
      -- CP-element group 93: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_305_Update/ca
      -- 
    ca_727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_305_inst_ack_1, ack => convTranspose_CP_39_elements(93)); -- 
    -- CP-element group 94:  transition  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	91 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (6) 
      -- CP-element group 94: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_313_sample_completed_
      -- CP-element group 94: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_313_update_start_
      -- CP-element group 94: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_313_Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_313_Sample/ra
      -- CP-element group 94: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_313_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_313_Update/cr
      -- 
    ra_736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_313_inst_ack_0, ack => convTranspose_CP_39_elements(94)); -- 
    cr_740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(94), ack => RPIPE_ConvTranspose_input_pipe_313_inst_req_1); -- 
    -- CP-element group 95:  fork  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95: 	98 
    -- CP-element group 95:  members (9) 
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_317_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_317_Sample/rr
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_326_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_326_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_326_Sample/rr
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_313_update_completed_
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_313_Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_313_Update/ca
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_317_sample_start_
      -- 
    ca_741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_313_inst_ack_1, ack => convTranspose_CP_39_elements(95)); -- 
    rr_749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(95), ack => type_cast_317_inst_req_0); -- 
    rr_763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(95), ack => RPIPE_ConvTranspose_input_pipe_326_inst_req_0); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_317_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_317_Sample/ra
      -- CP-element group 96: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_317_sample_completed_
      -- 
    ra_750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_317_inst_ack_0, ack => convTranspose_CP_39_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	0 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	118 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_317_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_317_Update/ca
      -- CP-element group 97: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_317_update_completed_
      -- 
    ca_755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_317_inst_ack_1, ack => convTranspose_CP_39_elements(97)); -- 
    -- CP-element group 98:  transition  input  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	95 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (6) 
      -- CP-element group 98: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_326_sample_completed_
      -- CP-element group 98: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_326_update_start_
      -- CP-element group 98: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_326_Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_326_Sample/ra
      -- CP-element group 98: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_326_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_326_Update/cr
      -- 
    ra_764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_326_inst_ack_0, ack => convTranspose_CP_39_elements(98)); -- 
    cr_768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(98), ack => RPIPE_ConvTranspose_input_pipe_326_inst_req_1); -- 
    -- CP-element group 99:  fork  transition  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: 	102 
    -- CP-element group 99:  members (9) 
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_326_update_completed_
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_326_Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_326_Update/ca
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_330_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_330_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_330_Sample/rr
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_338_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_338_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_338_Sample/rr
      -- 
    ca_769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_326_inst_ack_1, ack => convTranspose_CP_39_elements(99)); -- 
    rr_777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(99), ack => type_cast_330_inst_req_0); -- 
    rr_791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(99), ack => RPIPE_ConvTranspose_input_pipe_338_inst_req_0); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_330_sample_completed_
      -- CP-element group 100: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_330_Sample/$exit
      -- CP-element group 100: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_330_Sample/ra
      -- 
    ra_778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_330_inst_ack_0, ack => convTranspose_CP_39_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	0 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	118 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_330_update_completed_
      -- CP-element group 101: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_330_Update/$exit
      -- CP-element group 101: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_330_Update/ca
      -- 
    ca_783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_330_inst_ack_1, ack => convTranspose_CP_39_elements(101)); -- 
    -- CP-element group 102:  transition  input  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	99 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102:  members (6) 
      -- CP-element group 102: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_338_sample_completed_
      -- CP-element group 102: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_338_update_start_
      -- CP-element group 102: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_338_Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_338_Sample/ra
      -- CP-element group 102: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_338_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_338_Update/cr
      -- 
    ra_792_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_338_inst_ack_0, ack => convTranspose_CP_39_elements(102)); -- 
    cr_796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(102), ack => RPIPE_ConvTranspose_input_pipe_338_inst_req_1); -- 
    -- CP-element group 103:  fork  transition  input  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103: 	106 
    -- CP-element group 103:  members (9) 
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_338_update_completed_
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_338_Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_338_Update/ca
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_342_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_342_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_342_Sample/rr
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_351_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_351_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_351_Sample/rr
      -- 
    ca_797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_338_inst_ack_1, ack => convTranspose_CP_39_elements(103)); -- 
    rr_805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(103), ack => type_cast_342_inst_req_0); -- 
    rr_819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(103), ack => RPIPE_ConvTranspose_input_pipe_351_inst_req_0); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_342_sample_completed_
      -- CP-element group 104: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_342_Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_342_Sample/ra
      -- 
    ra_806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_342_inst_ack_0, ack => convTranspose_CP_39_elements(104)); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	0 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	118 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_342_update_completed_
      -- CP-element group 105: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_342_Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_342_Update/ca
      -- 
    ca_811_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_342_inst_ack_1, ack => convTranspose_CP_39_elements(105)); -- 
    -- CP-element group 106:  transition  input  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	103 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (6) 
      -- CP-element group 106: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_351_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_351_update_start_
      -- CP-element group 106: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_351_Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_351_Sample/ra
      -- CP-element group 106: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_351_Update/$entry
      -- CP-element group 106: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_351_Update/cr
      -- 
    ra_820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_351_inst_ack_0, ack => convTranspose_CP_39_elements(106)); -- 
    cr_824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(106), ack => RPIPE_ConvTranspose_input_pipe_351_inst_req_1); -- 
    -- CP-element group 107:  fork  transition  input  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107: 	110 
    -- CP-element group 107:  members (9) 
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_351_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_351_Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_351_Update/ca
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_355_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_355_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_355_Sample/rr
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_363_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_363_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_363_Sample/rr
      -- 
    ca_825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_351_inst_ack_1, ack => convTranspose_CP_39_elements(107)); -- 
    rr_833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(107), ack => type_cast_355_inst_req_0); -- 
    rr_847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(107), ack => RPIPE_ConvTranspose_input_pipe_363_inst_req_0); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_355_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_355_Sample/$exit
      -- CP-element group 108: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_355_Sample/ra
      -- 
    ra_834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_355_inst_ack_0, ack => convTranspose_CP_39_elements(108)); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	0 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	118 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_355_update_completed_
      -- CP-element group 109: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_355_Update/$exit
      -- CP-element group 109: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_355_Update/ca
      -- 
    ca_839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_355_inst_ack_1, ack => convTranspose_CP_39_elements(109)); -- 
    -- CP-element group 110:  transition  input  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	107 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (6) 
      -- CP-element group 110: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_363_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_363_update_start_
      -- CP-element group 110: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_363_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_363_Sample/ra
      -- CP-element group 110: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_363_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_363_Update/cr
      -- 
    ra_848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_363_inst_ack_0, ack => convTranspose_CP_39_elements(110)); -- 
    cr_852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(110), ack => RPIPE_ConvTranspose_input_pipe_363_inst_req_1); -- 
    -- CP-element group 111:  fork  transition  input  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111: 	114 
    -- CP-element group 111:  members (9) 
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_363_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_363_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_363_Update/ca
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_367_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_367_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_367_Sample/rr
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_376_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_376_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_376_Sample/rr
      -- 
    ca_853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_363_inst_ack_1, ack => convTranspose_CP_39_elements(111)); -- 
    rr_861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(111), ack => type_cast_367_inst_req_0); -- 
    rr_875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(111), ack => RPIPE_ConvTranspose_input_pipe_376_inst_req_0); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_367_sample_completed_
      -- CP-element group 112: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_367_Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_367_Sample/ra
      -- 
    ra_862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_367_inst_ack_0, ack => convTranspose_CP_39_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	0 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	118 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_367_update_completed_
      -- CP-element group 113: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_367_Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_367_Update/ca
      -- 
    ca_867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_367_inst_ack_1, ack => convTranspose_CP_39_elements(113)); -- 
    -- CP-element group 114:  transition  input  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	111 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (6) 
      -- CP-element group 114: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_376_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_376_update_start_
      -- CP-element group 114: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_376_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_376_Sample/ra
      -- CP-element group 114: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_376_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_376_Update/cr
      -- 
    ra_876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_376_inst_ack_0, ack => convTranspose_CP_39_elements(114)); -- 
    cr_880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(114), ack => RPIPE_ConvTranspose_input_pipe_376_inst_req_1); -- 
    -- CP-element group 115:  transition  input  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (6) 
      -- CP-element group 115: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_376_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_376_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_376_Update/ca
      -- CP-element group 115: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_380_sample_start_
      -- CP-element group 115: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_380_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_380_Sample/rr
      -- 
    ca_881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_376_inst_ack_1, ack => convTranspose_CP_39_elements(115)); -- 
    rr_889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(115), ack => type_cast_380_inst_req_0); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_380_sample_completed_
      -- CP-element group 116: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_380_Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_380_Sample/ra
      -- 
    ra_890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_380_inst_ack_0, ack => convTranspose_CP_39_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	0 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_380_update_completed_
      -- CP-element group 117: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_380_Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_380_Update/ca
      -- 
    ca_895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_380_inst_ack_1, ack => convTranspose_CP_39_elements(117)); -- 
    -- CP-element group 118:  branch  join  transition  place  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	68 
    -- CP-element group 118: 	62 
    -- CP-element group 118: 	65 
    -- CP-element group 118: 	59 
    -- CP-element group 118: 	71 
    -- CP-element group 118: 	74 
    -- CP-element group 118: 	77 
    -- CP-element group 118: 	81 
    -- CP-element group 118: 	85 
    -- CP-element group 118: 	89 
    -- CP-element group 118: 	93 
    -- CP-element group 118: 	97 
    -- CP-element group 118: 	101 
    -- CP-element group 118: 	105 
    -- CP-element group 118: 	109 
    -- CP-element group 118: 	113 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118: 	120 
    -- CP-element group 118:  members (10) 
      -- CP-element group 118: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393__exit__
      -- CP-element group 118: 	 branch_block_stmt_33/if_stmt_394__entry__
      -- CP-element group 118: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/$exit
      -- CP-element group 118: 	 branch_block_stmt_33/if_stmt_394_dead_link/$entry
      -- CP-element group 118: 	 branch_block_stmt_33/if_stmt_394_eval_test/$entry
      -- CP-element group 118: 	 branch_block_stmt_33/if_stmt_394_eval_test/$exit
      -- CP-element group 118: 	 branch_block_stmt_33/if_stmt_394_eval_test/branch_req
      -- CP-element group 118: 	 branch_block_stmt_33/R_cmp417_395_place
      -- CP-element group 118: 	 branch_block_stmt_33/if_stmt_394_if_link/$entry
      -- CP-element group 118: 	 branch_block_stmt_33/if_stmt_394_else_link/$entry
      -- 
    branch_req_903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(118), ack => if_stmt_394_branch_req_0); -- 
    convTranspose_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(68) & convTranspose_CP_39_elements(62) & convTranspose_CP_39_elements(65) & convTranspose_CP_39_elements(59) & convTranspose_CP_39_elements(71) & convTranspose_CP_39_elements(74) & convTranspose_CP_39_elements(77) & convTranspose_CP_39_elements(81) & convTranspose_CP_39_elements(85) & convTranspose_CP_39_elements(89) & convTranspose_CP_39_elements(93) & convTranspose_CP_39_elements(97) & convTranspose_CP_39_elements(101) & convTranspose_CP_39_elements(105) & convTranspose_CP_39_elements(109) & convTranspose_CP_39_elements(113) & convTranspose_CP_39_elements(117);
      gj_convTranspose_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	123 
    -- CP-element group 119: 	124 
    -- CP-element group 119:  members (18) 
      -- CP-element group 119: 	 branch_block_stmt_33/merge_stmt_415__exit__
      -- CP-element group 119: 	 branch_block_stmt_33/assign_stmt_421_to_assign_stmt_450__entry__
      -- CP-element group 119: 	 branch_block_stmt_33/if_stmt_394_if_link/$exit
      -- CP-element group 119: 	 branch_block_stmt_33/if_stmt_394_if_link/if_choice_transition
      -- CP-element group 119: 	 branch_block_stmt_33/entry_bbx_xnph419
      -- CP-element group 119: 	 branch_block_stmt_33/assign_stmt_421_to_assign_stmt_450/$entry
      -- CP-element group 119: 	 branch_block_stmt_33/assign_stmt_421_to_assign_stmt_450/type_cast_436_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_33/assign_stmt_421_to_assign_stmt_450/type_cast_436_update_start_
      -- CP-element group 119: 	 branch_block_stmt_33/assign_stmt_421_to_assign_stmt_450/type_cast_436_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_33/assign_stmt_421_to_assign_stmt_450/type_cast_436_Sample/rr
      -- CP-element group 119: 	 branch_block_stmt_33/assign_stmt_421_to_assign_stmt_450/type_cast_436_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_33/assign_stmt_421_to_assign_stmt_450/type_cast_436_Update/cr
      -- CP-element group 119: 	 branch_block_stmt_33/merge_stmt_415_PhiReqMerge
      -- CP-element group 119: 	 branch_block_stmt_33/merge_stmt_415_PhiAck/dummy
      -- CP-element group 119: 	 branch_block_stmt_33/merge_stmt_415_PhiAck/$exit
      -- CP-element group 119: 	 branch_block_stmt_33/merge_stmt_415_PhiAck/$entry
      -- CP-element group 119: 	 branch_block_stmt_33/entry_bbx_xnph419_PhiReq/$exit
      -- CP-element group 119: 	 branch_block_stmt_33/entry_bbx_xnph419_PhiReq/$entry
      -- 
    if_choice_transition_908_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_394_branch_ack_1, ack => convTranspose_CP_39_elements(119)); -- 
    rr_947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(119), ack => type_cast_436_inst_req_0); -- 
    cr_952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(119), ack => type_cast_436_inst_req_1); -- 
    -- CP-element group 120:  transition  place  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	118 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	398 
    -- CP-element group 120:  members (5) 
      -- CP-element group 120: 	 branch_block_stmt_33/if_stmt_394_else_link/$exit
      -- CP-element group 120: 	 branch_block_stmt_33/if_stmt_394_else_link/else_choice_transition
      -- CP-element group 120: 	 branch_block_stmt_33/entry_forx_xcond176x_xpreheader
      -- CP-element group 120: 	 branch_block_stmt_33/entry_forx_xcond176x_xpreheader_PhiReq/$exit
      -- CP-element group 120: 	 branch_block_stmt_33/entry_forx_xcond176x_xpreheader_PhiReq/$entry
      -- 
    else_choice_transition_912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_394_branch_ack_0, ack => convTranspose_CP_39_elements(120)); -- 
    -- CP-element group 121:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	398 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	167 
    -- CP-element group 121: 	168 
    -- CP-element group 121:  members (18) 
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_628_to_assign_stmt_657/type_cast_643_Sample/$entry
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_628_to_assign_stmt_657/type_cast_643_Sample/rr
      -- CP-element group 121: 	 branch_block_stmt_33/merge_stmt_622__exit__
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_628_to_assign_stmt_657__entry__
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_628_to_assign_stmt_657/type_cast_643_update_start_
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_628_to_assign_stmt_657/type_cast_643_Update/cr
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_628_to_assign_stmt_657/type_cast_643_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_628_to_assign_stmt_657/$entry
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_628_to_assign_stmt_657/type_cast_643_Update/$entry
      -- CP-element group 121: 	 branch_block_stmt_33/merge_stmt_622_PhiReqMerge
      -- CP-element group 121: 	 branch_block_stmt_33/if_stmt_409_if_link/$exit
      -- CP-element group 121: 	 branch_block_stmt_33/if_stmt_409_if_link/if_choice_transition
      -- CP-element group 121: 	 branch_block_stmt_33/forx_xcond176x_xpreheader_bbx_xnph415
      -- CP-element group 121: 	 branch_block_stmt_33/forx_xcond176x_xpreheader_bbx_xnph415_PhiReq/$entry
      -- CP-element group 121: 	 branch_block_stmt_33/forx_xcond176x_xpreheader_bbx_xnph415_PhiReq/$exit
      -- CP-element group 121: 	 branch_block_stmt_33/merge_stmt_622_PhiAck/$entry
      -- CP-element group 121: 	 branch_block_stmt_33/merge_stmt_622_PhiAck/$exit
      -- CP-element group 121: 	 branch_block_stmt_33/merge_stmt_622_PhiAck/dummy
      -- 
    if_choice_transition_930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_409_branch_ack_1, ack => convTranspose_CP_39_elements(121)); -- 
    rr_1306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(121), ack => type_cast_643_inst_req_0); -- 
    cr_1311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(121), ack => type_cast_643_inst_req_1); -- 
    -- CP-element group 122:  transition  place  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	398 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	411 
    -- CP-element group 122:  members (5) 
      -- CP-element group 122: 	 branch_block_stmt_33/if_stmt_409_else_link/$exit
      -- CP-element group 122: 	 branch_block_stmt_33/if_stmt_409_else_link/else_choice_transition
      -- CP-element group 122: 	 branch_block_stmt_33/forx_xcond176x_xpreheader_forx_xend236
      -- CP-element group 122: 	 branch_block_stmt_33/forx_xcond176x_xpreheader_forx_xend236_PhiReq/$exit
      -- CP-element group 122: 	 branch_block_stmt_33/forx_xcond176x_xpreheader_forx_xend236_PhiReq/$entry
      -- 
    else_choice_transition_934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_409_branch_ack_0, ack => convTranspose_CP_39_elements(122)); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	119 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_33/assign_stmt_421_to_assign_stmt_450/type_cast_436_sample_completed_
      -- CP-element group 123: 	 branch_block_stmt_33/assign_stmt_421_to_assign_stmt_450/type_cast_436_Sample/$exit
      -- CP-element group 123: 	 branch_block_stmt_33/assign_stmt_421_to_assign_stmt_450/type_cast_436_Sample/ra
      -- 
    ra_948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_436_inst_ack_0, ack => convTranspose_CP_39_elements(123)); -- 
    -- CP-element group 124:  transition  place  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	119 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	399 
    -- CP-element group 124:  members (9) 
      -- CP-element group 124: 	 branch_block_stmt_33/assign_stmt_421_to_assign_stmt_450__exit__
      -- CP-element group 124: 	 branch_block_stmt_33/bbx_xnph419_forx_xbody
      -- CP-element group 124: 	 branch_block_stmt_33/assign_stmt_421_to_assign_stmt_450/$exit
      -- CP-element group 124: 	 branch_block_stmt_33/assign_stmt_421_to_assign_stmt_450/type_cast_436_update_completed_
      -- CP-element group 124: 	 branch_block_stmt_33/assign_stmt_421_to_assign_stmt_450/type_cast_436_Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_33/assign_stmt_421_to_assign_stmt_450/type_cast_436_Update/ca
      -- CP-element group 124: 	 branch_block_stmt_33/bbx_xnph419_forx_xbody_PhiReq/phi_stmt_453/phi_stmt_453_sources/$entry
      -- CP-element group 124: 	 branch_block_stmt_33/bbx_xnph419_forx_xbody_PhiReq/phi_stmt_453/$entry
      -- CP-element group 124: 	 branch_block_stmt_33/bbx_xnph419_forx_xbody_PhiReq/$entry
      -- 
    ca_953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_436_inst_ack_1, ack => convTranspose_CP_39_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	404 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	164 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_final_index_sum_regn_sample_complete
      -- CP-element group 125: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_final_index_sum_regn_Sample/$exit
      -- CP-element group 125: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_final_index_sum_regn_Sample/ack
      -- 
    ack_982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_465_index_offset_ack_0, ack => convTranspose_CP_39_elements(125)); -- 
    -- CP-element group 126:  transition  input  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	404 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (11) 
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/addr_of_466_sample_start_
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_root_address_calculated
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_offset_calculated
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_final_index_sum_regn_Update/$exit
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_final_index_sum_regn_Update/ack
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_base_plus_offset/$entry
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_base_plus_offset/$exit
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_base_plus_offset/sum_rename_req
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_base_plus_offset/sum_rename_ack
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/addr_of_466_request/$entry
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/addr_of_466_request/req
      -- 
    ack_987_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_465_index_offset_ack_1, ack => convTranspose_CP_39_elements(126)); -- 
    req_996_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_996_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(126), ack => addr_of_466_final_reg_req_0); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/addr_of_466_sample_completed_
      -- CP-element group 127: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/addr_of_466_request/$exit
      -- CP-element group 127: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/addr_of_466_request/ack
      -- 
    ack_997_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_466_final_reg_ack_0, ack => convTranspose_CP_39_elements(127)); -- 
    -- CP-element group 128:  fork  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	404 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	161 
    -- CP-element group 128:  members (19) 
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_word_addrgen/root_register_ack
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_word_addrgen/root_register_req
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_word_addrgen/$exit
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_word_addrgen/$entry
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_base_plus_offset/sum_rename_ack
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_base_plus_offset/sum_rename_req
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_base_plus_offset/$exit
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_base_plus_offset/$entry
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_base_addr_resize/base_resize_ack
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_base_addr_resize/base_resize_req
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_base_addr_resize/$exit
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_base_addr_resize/$entry
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_base_address_resized
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_root_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_word_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_base_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/addr_of_466_update_completed_
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/addr_of_466_complete/$exit
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/addr_of_466_complete/ack
      -- 
    ack_1002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_466_final_reg_ack_1, ack => convTranspose_CP_39_elements(128)); -- 
    -- CP-element group 129:  transition  input  output  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	404 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (6) 
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_469_sample_completed_
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_469_update_start_
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_469_Sample/$exit
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_469_Sample/ra
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_469_Update/$entry
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_469_Update/cr
      -- 
    ra_1011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_469_inst_ack_0, ack => convTranspose_CP_39_elements(129)); -- 
    cr_1015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(129), ack => RPIPE_ConvTranspose_input_pipe_469_inst_req_1); -- 
    -- CP-element group 130:  fork  transition  input  output  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130: 	133 
    -- CP-element group 130:  members (9) 
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_469_update_completed_
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_469_Update/$exit
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_469_Update/ca
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_473_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_473_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_473_Sample/rr
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_482_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_482_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_482_Sample/rr
      -- 
    ca_1016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_469_inst_ack_1, ack => convTranspose_CP_39_elements(130)); -- 
    rr_1024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(130), ack => type_cast_473_inst_req_0); -- 
    rr_1038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(130), ack => RPIPE_ConvTranspose_input_pipe_482_inst_req_0); -- 
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_473_sample_completed_
      -- CP-element group 131: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_473_Sample/$exit
      -- CP-element group 131: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_473_Sample/ra
      -- 
    ra_1025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_473_inst_ack_0, ack => convTranspose_CP_39_elements(131)); -- 
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	404 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	161 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_473_update_completed_
      -- CP-element group 132: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_473_Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_473_Update/ca
      -- 
    ca_1030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_473_inst_ack_1, ack => convTranspose_CP_39_elements(132)); -- 
    -- CP-element group 133:  transition  input  output  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	130 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133:  members (6) 
      -- CP-element group 133: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_482_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_482_update_start_
      -- CP-element group 133: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_482_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_482_Sample/ra
      -- CP-element group 133: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_482_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_482_Update/cr
      -- 
    ra_1039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_482_inst_ack_0, ack => convTranspose_CP_39_elements(133)); -- 
    cr_1043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(133), ack => RPIPE_ConvTranspose_input_pipe_482_inst_req_1); -- 
    -- CP-element group 134:  fork  transition  input  output  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134: 	137 
    -- CP-element group 134:  members (9) 
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_482_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_482_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_482_Update/ca
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_486_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_486_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_486_Sample/rr
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_500_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_500_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_500_Sample/rr
      -- 
    ca_1044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_482_inst_ack_1, ack => convTranspose_CP_39_elements(134)); -- 
    rr_1052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(134), ack => type_cast_486_inst_req_0); -- 
    rr_1066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(134), ack => RPIPE_ConvTranspose_input_pipe_500_inst_req_0); -- 
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	134 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_486_sample_completed_
      -- CP-element group 135: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_486_Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_486_Sample/ra
      -- 
    ra_1053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_486_inst_ack_0, ack => convTranspose_CP_39_elements(135)); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	404 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	161 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_486_update_completed_
      -- CP-element group 136: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_486_Update/$exit
      -- CP-element group 136: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_486_Update/ca
      -- 
    ca_1058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_486_inst_ack_1, ack => convTranspose_CP_39_elements(136)); -- 
    -- CP-element group 137:  transition  input  output  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	134 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137:  members (6) 
      -- CP-element group 137: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_500_sample_completed_
      -- CP-element group 137: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_500_update_start_
      -- CP-element group 137: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_500_Sample/$exit
      -- CP-element group 137: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_500_Sample/ra
      -- CP-element group 137: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_500_Update/$entry
      -- CP-element group 137: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_500_Update/cr
      -- 
    ra_1067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_500_inst_ack_0, ack => convTranspose_CP_39_elements(137)); -- 
    cr_1071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(137), ack => RPIPE_ConvTranspose_input_pipe_500_inst_req_1); -- 
    -- CP-element group 138:  fork  transition  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	139 
    -- CP-element group 138: 	141 
    -- CP-element group 138:  members (9) 
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_518_Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_518_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_518_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_500_update_completed_
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_500_Update/$exit
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_500_Update/ca
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_504_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_504_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_504_Sample/rr
      -- 
    ca_1072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_500_inst_ack_1, ack => convTranspose_CP_39_elements(138)); -- 
    rr_1080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(138), ack => type_cast_504_inst_req_0); -- 
    rr_1094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(138), ack => RPIPE_ConvTranspose_input_pipe_518_inst_req_0); -- 
    -- CP-element group 139:  transition  input  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	138 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_504_Sample/ra
      -- CP-element group 139: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_504_sample_completed_
      -- CP-element group 139: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_504_Sample/$exit
      -- 
    ra_1081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_504_inst_ack_0, ack => convTranspose_CP_39_elements(139)); -- 
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	404 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	161 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_504_Update/ca
      -- CP-element group 140: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_504_Update/$exit
      -- CP-element group 140: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_504_update_completed_
      -- 
    ca_1086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_504_inst_ack_1, ack => convTranspose_CP_39_elements(140)); -- 
    -- CP-element group 141:  transition  input  output  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	138 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	142 
    -- CP-element group 141:  members (6) 
      -- CP-element group 141: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_518_update_start_
      -- CP-element group 141: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_518_Sample/$exit
      -- CP-element group 141: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_518_Update/cr
      -- CP-element group 141: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_518_Update/$entry
      -- CP-element group 141: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_518_Sample/ra
      -- CP-element group 141: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_518_sample_completed_
      -- 
    ra_1095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_518_inst_ack_0, ack => convTranspose_CP_39_elements(141)); -- 
    cr_1099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(141), ack => RPIPE_ConvTranspose_input_pipe_518_inst_req_1); -- 
    -- CP-element group 142:  fork  transition  input  output  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	141 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	143 
    -- CP-element group 142: 	145 
    -- CP-element group 142:  members (9) 
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_522_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_518_Update/ca
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_518_Update/$exit
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_536_Sample/rr
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_536_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_536_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_522_Sample/rr
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_522_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_518_update_completed_
      -- 
    ca_1100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_518_inst_ack_1, ack => convTranspose_CP_39_elements(142)); -- 
    rr_1108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(142), ack => type_cast_522_inst_req_0); -- 
    rr_1122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(142), ack => RPIPE_ConvTranspose_input_pipe_536_inst_req_0); -- 
    -- CP-element group 143:  transition  input  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	142 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_522_sample_completed_
      -- CP-element group 143: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_522_Sample/ra
      -- CP-element group 143: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_522_Sample/$exit
      -- 
    ra_1109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_522_inst_ack_0, ack => convTranspose_CP_39_elements(143)); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	404 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	161 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_522_update_completed_
      -- CP-element group 144: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_522_Update/ca
      -- CP-element group 144: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_522_Update/$exit
      -- 
    ca_1114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_522_inst_ack_1, ack => convTranspose_CP_39_elements(144)); -- 
    -- CP-element group 145:  transition  input  output  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	142 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145:  members (6) 
      -- CP-element group 145: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_536_Update/cr
      -- CP-element group 145: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_536_Update/$entry
      -- CP-element group 145: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_536_Sample/ra
      -- CP-element group 145: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_536_Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_536_update_start_
      -- CP-element group 145: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_536_sample_completed_
      -- 
    ra_1123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_536_inst_ack_0, ack => convTranspose_CP_39_elements(145)); -- 
    cr_1127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(145), ack => RPIPE_ConvTranspose_input_pipe_536_inst_req_1); -- 
    -- CP-element group 146:  fork  transition  input  output  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	145 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	147 
    -- CP-element group 146: 	149 
    -- CP-element group 146:  members (9) 
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_554_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_554_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_554_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_540_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_540_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_540_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_536_Update/ca
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_536_Update/$exit
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_536_update_completed_
      -- 
    ca_1128_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_536_inst_ack_1, ack => convTranspose_CP_39_elements(146)); -- 
    rr_1136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(146), ack => type_cast_540_inst_req_0); -- 
    rr_1150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(146), ack => RPIPE_ConvTranspose_input_pipe_554_inst_req_0); -- 
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	146 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_540_Sample/ra
      -- CP-element group 147: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_540_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_540_sample_completed_
      -- 
    ra_1137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_540_inst_ack_0, ack => convTranspose_CP_39_elements(147)); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	404 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	161 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_540_Update/ca
      -- CP-element group 148: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_540_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_540_update_completed_
      -- 
    ca_1142_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_540_inst_ack_1, ack => convTranspose_CP_39_elements(148)); -- 
    -- CP-element group 149:  transition  input  output  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	146 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	150 
    -- CP-element group 149:  members (6) 
      -- CP-element group 149: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_554_Sample/ra
      -- CP-element group 149: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_554_Update/cr
      -- CP-element group 149: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_554_Update/$entry
      -- CP-element group 149: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_554_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_554_update_start_
      -- CP-element group 149: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_554_sample_completed_
      -- 
    ra_1151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_554_inst_ack_0, ack => convTranspose_CP_39_elements(149)); -- 
    cr_1155_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1155_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(149), ack => RPIPE_ConvTranspose_input_pipe_554_inst_req_1); -- 
    -- CP-element group 150:  fork  transition  input  output  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	149 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	151 
    -- CP-element group 150: 	153 
    -- CP-element group 150:  members (9) 
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_572_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_572_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_572_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_558_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_558_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_558_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_554_Update/ca
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_554_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_554_update_completed_
      -- 
    ca_1156_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_554_inst_ack_1, ack => convTranspose_CP_39_elements(150)); -- 
    rr_1164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(150), ack => type_cast_558_inst_req_0); -- 
    rr_1178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(150), ack => RPIPE_ConvTranspose_input_pipe_572_inst_req_0); -- 
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	150 
    -- CP-element group 151: successors 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_558_Sample/ra
      -- CP-element group 151: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_558_sample_completed_
      -- CP-element group 151: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_558_Sample/$exit
      -- 
    ra_1165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_558_inst_ack_0, ack => convTranspose_CP_39_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	404 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	161 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_558_Update/ca
      -- CP-element group 152: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_558_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_558_update_completed_
      -- 
    ca_1170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_558_inst_ack_1, ack => convTranspose_CP_39_elements(152)); -- 
    -- CP-element group 153:  transition  input  output  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	150 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153:  members (6) 
      -- CP-element group 153: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_572_sample_completed_
      -- CP-element group 153: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_572_Update/cr
      -- CP-element group 153: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_572_Update/$entry
      -- CP-element group 153: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_572_Sample/ra
      -- CP-element group 153: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_572_Sample/$exit
      -- CP-element group 153: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_572_update_start_
      -- 
    ra_1179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_572_inst_ack_0, ack => convTranspose_CP_39_elements(153)); -- 
    cr_1183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(153), ack => RPIPE_ConvTranspose_input_pipe_572_inst_req_1); -- 
    -- CP-element group 154:  fork  transition  input  output  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154: 	157 
    -- CP-element group 154:  members (9) 
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_576_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_572_Update/ca
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_572_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_572_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_590_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_590_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_590_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_576_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_576_Sample/$entry
      -- 
    ca_1184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_572_inst_ack_1, ack => convTranspose_CP_39_elements(154)); -- 
    rr_1192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(154), ack => type_cast_576_inst_req_0); -- 
    rr_1206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(154), ack => RPIPE_ConvTranspose_input_pipe_590_inst_req_0); -- 
    -- CP-element group 155:  transition  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_576_Sample/ra
      -- CP-element group 155: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_576_Sample/$exit
      -- CP-element group 155: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_576_sample_completed_
      -- 
    ra_1193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_576_inst_ack_0, ack => convTranspose_CP_39_elements(155)); -- 
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	404 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	161 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_576_Update/ca
      -- CP-element group 156: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_576_Update/$exit
      -- CP-element group 156: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_576_update_completed_
      -- 
    ca_1198_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_576_inst_ack_1, ack => convTranspose_CP_39_elements(156)); -- 
    -- CP-element group 157:  transition  input  output  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	154 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	158 
    -- CP-element group 157:  members (6) 
      -- CP-element group 157: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_590_Update/cr
      -- CP-element group 157: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_590_Update/$entry
      -- CP-element group 157: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_590_Sample/ra
      -- CP-element group 157: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_590_Sample/$exit
      -- CP-element group 157: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_590_update_start_
      -- CP-element group 157: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_590_sample_completed_
      -- 
    ra_1207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_590_inst_ack_0, ack => convTranspose_CP_39_elements(157)); -- 
    cr_1211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(157), ack => RPIPE_ConvTranspose_input_pipe_590_inst_req_1); -- 
    -- CP-element group 158:  transition  input  output  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	157 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	159 
    -- CP-element group 158:  members (6) 
      -- CP-element group 158: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_594_Sample/$entry
      -- CP-element group 158: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_594_Sample/rr
      -- CP-element group 158: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_594_sample_start_
      -- CP-element group 158: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_590_Update/ca
      -- CP-element group 158: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_590_Update/$exit
      -- CP-element group 158: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_590_update_completed_
      -- 
    ca_1212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_590_inst_ack_1, ack => convTranspose_CP_39_elements(158)); -- 
    rr_1220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(158), ack => type_cast_594_inst_req_0); -- 
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	158 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_594_Sample/$exit
      -- CP-element group 159: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_594_sample_completed_
      -- CP-element group 159: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_594_Sample/ra
      -- 
    ra_1221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_594_inst_ack_0, ack => convTranspose_CP_39_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	404 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	161 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_594_update_completed_
      -- CP-element group 160: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_594_Update/ca
      -- CP-element group 160: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_594_Update/$exit
      -- 
    ca_1226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_594_inst_ack_1, ack => convTranspose_CP_39_elements(160)); -- 
    -- CP-element group 161:  join  transition  output  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	128 
    -- CP-element group 161: 	132 
    -- CP-element group 161: 	136 
    -- CP-element group 161: 	140 
    -- CP-element group 161: 	144 
    -- CP-element group 161: 	148 
    -- CP-element group 161: 	152 
    -- CP-element group 161: 	156 
    -- CP-element group 161: 	160 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161:  members (9) 
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_Sample/word_access_start/word_0/rr
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_Sample/word_access_start/word_0/$entry
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_Sample/word_access_start/$entry
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_Sample/ptr_deref_602_Split/split_ack
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_Sample/ptr_deref_602_Split/split_req
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_Sample/ptr_deref_602_Split/$exit
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_Sample/ptr_deref_602_Split/$entry
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_Sample/$entry
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_sample_start_
      -- 
    rr_1264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(161), ack => ptr_deref_602_store_0_req_0); -- 
    convTranspose_cp_element_group_161: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_161"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(128) & convTranspose_CP_39_elements(132) & convTranspose_CP_39_elements(136) & convTranspose_CP_39_elements(140) & convTranspose_CP_39_elements(144) & convTranspose_CP_39_elements(148) & convTranspose_CP_39_elements(152) & convTranspose_CP_39_elements(156) & convTranspose_CP_39_elements(160);
      gj_convTranspose_cp_element_group_161 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(161), clk => clk, reset => reset); --
    end block;
    -- CP-element group 162:  transition  input  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	161 
    -- CP-element group 162: successors 
    -- CP-element group 162:  members (5) 
      -- CP-element group 162: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_Sample/word_access_start/word_0/ra
      -- CP-element group 162: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_Sample/word_access_start/word_0/$exit
      -- CP-element group 162: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_Sample/word_access_start/$exit
      -- CP-element group 162: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_Sample/$exit
      -- CP-element group 162: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_sample_completed_
      -- 
    ra_1265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_602_store_0_ack_0, ack => convTranspose_CP_39_elements(162)); -- 
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	404 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	164 
    -- CP-element group 163:  members (5) 
      -- CP-element group 163: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_Update/$exit
      -- CP-element group 163: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_update_completed_
      -- CP-element group 163: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_Update/word_access_complete/word_0/ca
      -- CP-element group 163: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_Update/word_access_complete/word_0/$exit
      -- CP-element group 163: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_Update/word_access_complete/$exit
      -- 
    ca_1276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_602_store_0_ack_1, ack => convTranspose_CP_39_elements(163)); -- 
    -- CP-element group 164:  branch  join  transition  place  output  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	163 
    -- CP-element group 164: 	125 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	165 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (10) 
      -- CP-element group 164: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615__exit__
      -- CP-element group 164: 	 branch_block_stmt_33/if_stmt_616__entry__
      -- CP-element group 164: 	 branch_block_stmt_33/if_stmt_616_else_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_33/if_stmt_616_if_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_33/R_exitcond3_617_place
      -- CP-element group 164: 	 branch_block_stmt_33/if_stmt_616_eval_test/branch_req
      -- CP-element group 164: 	 branch_block_stmt_33/if_stmt_616_eval_test/$exit
      -- CP-element group 164: 	 branch_block_stmt_33/if_stmt_616_eval_test/$entry
      -- CP-element group 164: 	 branch_block_stmt_33/if_stmt_616_dead_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/$exit
      -- 
    branch_req_1284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(164), ack => if_stmt_616_branch_req_0); -- 
    convTranspose_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(163) & convTranspose_CP_39_elements(125);
      gj_convTranspose_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  merge  transition  place  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	164 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	398 
    -- CP-element group 165:  members (13) 
      -- CP-element group 165: 	 branch_block_stmt_33/merge_stmt_400__exit__
      -- CP-element group 165: 	 branch_block_stmt_33/forx_xcond176x_xpreheaderx_xloopexit_forx_xcond176x_xpreheader
      -- CP-element group 165: 	 branch_block_stmt_33/forx_xbody_forx_xcond176x_xpreheaderx_xloopexit
      -- CP-element group 165: 	 branch_block_stmt_33/merge_stmt_400_PhiReqMerge
      -- CP-element group 165: 	 branch_block_stmt_33/if_stmt_616_if_link/if_choice_transition
      -- CP-element group 165: 	 branch_block_stmt_33/if_stmt_616_if_link/$exit
      -- CP-element group 165: 	 branch_block_stmt_33/merge_stmt_400_PhiAck/$entry
      -- CP-element group 165: 	 branch_block_stmt_33/merge_stmt_400_PhiAck/$exit
      -- CP-element group 165: 	 branch_block_stmt_33/forx_xbody_forx_xcond176x_xpreheaderx_xloopexit_PhiReq/$entry
      -- CP-element group 165: 	 branch_block_stmt_33/merge_stmt_400_PhiAck/dummy
      -- CP-element group 165: 	 branch_block_stmt_33/forx_xbody_forx_xcond176x_xpreheaderx_xloopexit_PhiReq/$exit
      -- CP-element group 165: 	 branch_block_stmt_33/forx_xcond176x_xpreheaderx_xloopexit_forx_xcond176x_xpreheader_PhiReq/$exit
      -- CP-element group 165: 	 branch_block_stmt_33/forx_xcond176x_xpreheaderx_xloopexit_forx_xcond176x_xpreheader_PhiReq/$entry
      -- 
    if_choice_transition_1289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_616_branch_ack_1, ack => convTranspose_CP_39_elements(165)); -- 
    -- CP-element group 166:  fork  transition  place  input  output  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	400 
    -- CP-element group 166: 	401 
    -- CP-element group 166:  members (12) 
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody_forx_xbody
      -- CP-element group 166: 	 branch_block_stmt_33/if_stmt_616_else_link/else_choice_transition
      -- CP-element group 166: 	 branch_block_stmt_33/if_stmt_616_else_link/$exit
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_453/phi_stmt_453_sources/type_cast_459/SplitProtocol/Update/cr
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_453/phi_stmt_453_sources/type_cast_459/SplitProtocol/Update/$entry
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_453/phi_stmt_453_sources/type_cast_459/SplitProtocol/Sample/rr
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_453/phi_stmt_453_sources/type_cast_459/SplitProtocol/Sample/$entry
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_453/phi_stmt_453_sources/type_cast_459/SplitProtocol/$entry
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_453/phi_stmt_453_sources/type_cast_459/$entry
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_453/phi_stmt_453_sources/$entry
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_453/$entry
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/$entry
      -- 
    else_choice_transition_1293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_616_branch_ack_0, ack => convTranspose_CP_39_elements(166)); -- 
    cr_3105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(166), ack => type_cast_459_inst_req_1); -- 
    rr_3100_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3100_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(166), ack => type_cast_459_inst_req_0); -- 
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	121 
    -- CP-element group 167: successors 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_33/assign_stmt_628_to_assign_stmt_657/type_cast_643_Sample/ra
      -- CP-element group 167: 	 branch_block_stmt_33/assign_stmt_628_to_assign_stmt_657/type_cast_643_Sample/$exit
      -- CP-element group 167: 	 branch_block_stmt_33/assign_stmt_628_to_assign_stmt_657/type_cast_643_sample_completed_
      -- 
    ra_1307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_643_inst_ack_0, ack => convTranspose_CP_39_elements(167)); -- 
    -- CP-element group 168:  transition  place  input  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	121 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	405 
    -- CP-element group 168:  members (9) 
      -- CP-element group 168: 	 branch_block_stmt_33/assign_stmt_628_to_assign_stmt_657__exit__
      -- CP-element group 168: 	 branch_block_stmt_33/bbx_xnph415_forx_xbody182
      -- CP-element group 168: 	 branch_block_stmt_33/assign_stmt_628_to_assign_stmt_657/type_cast_643_Update/ca
      -- CP-element group 168: 	 branch_block_stmt_33/assign_stmt_628_to_assign_stmt_657/type_cast_643_update_completed_
      -- CP-element group 168: 	 branch_block_stmt_33/assign_stmt_628_to_assign_stmt_657/$exit
      -- CP-element group 168: 	 branch_block_stmt_33/assign_stmt_628_to_assign_stmt_657/type_cast_643_Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_33/bbx_xnph415_forx_xbody182_PhiReq/$entry
      -- CP-element group 168: 	 branch_block_stmt_33/bbx_xnph415_forx_xbody182_PhiReq/phi_stmt_660/$entry
      -- CP-element group 168: 	 branch_block_stmt_33/bbx_xnph415_forx_xbody182_PhiReq/phi_stmt_660/phi_stmt_660_sources/$entry
      -- 
    ca_1312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_643_inst_ack_1, ack => convTranspose_CP_39_elements(168)); -- 
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	410 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	208 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_final_index_sum_regn_sample_complete
      -- CP-element group 169: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_final_index_sum_regn_Sample/ack
      -- CP-element group 169: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_final_index_sum_regn_Sample/$exit
      -- 
    ack_1341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_672_index_offset_ack_0, ack => convTranspose_CP_39_elements(169)); -- 
    -- CP-element group 170:  transition  input  output  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	410 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	171 
    -- CP-element group 170:  members (11) 
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_base_plus_offset/$exit
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_base_plus_offset/$entry
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/addr_of_673_request/req
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_final_index_sum_regn_Update/ack
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/addr_of_673_request/$entry
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_final_index_sum_regn_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_base_plus_offset/sum_rename_ack
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_base_plus_offset/sum_rename_req
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_offset_calculated
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_root_address_calculated
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/addr_of_673_sample_start_
      -- 
    ack_1346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_672_index_offset_ack_1, ack => convTranspose_CP_39_elements(170)); -- 
    req_1355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(170), ack => addr_of_673_final_reg_req_0); -- 
    -- CP-element group 171:  transition  input  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	170 
    -- CP-element group 171: successors 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/addr_of_673_request/ack
      -- CP-element group 171: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/addr_of_673_request/$exit
      -- CP-element group 171: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/addr_of_673_sample_completed_
      -- 
    ack_1356_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_673_final_reg_ack_0, ack => convTranspose_CP_39_elements(171)); -- 
    -- CP-element group 172:  fork  transition  input  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	410 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	205 
    -- CP-element group 172:  members (19) 
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/addr_of_673_complete/$exit
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/addr_of_673_complete/ack
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/addr_of_673_update_completed_
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_base_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_word_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_root_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_base_address_resized
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_base_addr_resize/$entry
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_base_addr_resize/$exit
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_base_addr_resize/base_resize_req
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_base_addr_resize/base_resize_ack
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_base_plus_offset/$entry
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_base_plus_offset/$exit
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_base_plus_offset/sum_rename_req
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_base_plus_offset/sum_rename_ack
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_word_addrgen/$entry
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_word_addrgen/$exit
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_word_addrgen/root_register_req
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_word_addrgen/root_register_ack
      -- 
    ack_1361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_673_final_reg_ack_1, ack => convTranspose_CP_39_elements(172)); -- 
    -- CP-element group 173:  transition  input  output  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	410 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	174 
    -- CP-element group 173:  members (6) 
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_676_update_start_
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_676_sample_completed_
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_676_Update/cr
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_676_Update/$entry
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_676_Sample/ra
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_676_Sample/$exit
      -- 
    ra_1370_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_676_inst_ack_0, ack => convTranspose_CP_39_elements(173)); -- 
    cr_1374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(173), ack => RPIPE_ConvTranspose_input_pipe_676_inst_req_1); -- 
    -- CP-element group 174:  fork  transition  input  output  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	173 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	175 
    -- CP-element group 174: 	177 
    -- CP-element group 174:  members (9) 
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_689_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_689_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_680_Sample/rr
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_680_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_689_Sample/rr
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_680_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_676_Update/ca
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_676_Update/$exit
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_676_update_completed_
      -- 
    ca_1375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_676_inst_ack_1, ack => convTranspose_CP_39_elements(174)); -- 
    rr_1383_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1383_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(174), ack => type_cast_680_inst_req_0); -- 
    rr_1397_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1397_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(174), ack => RPIPE_ConvTranspose_input_pipe_689_inst_req_0); -- 
    -- CP-element group 175:  transition  input  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	174 
    -- CP-element group 175: successors 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_680_Sample/ra
      -- CP-element group 175: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_680_Sample/$exit
      -- CP-element group 175: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_680_sample_completed_
      -- 
    ra_1384_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_680_inst_ack_0, ack => convTranspose_CP_39_elements(175)); -- 
    -- CP-element group 176:  transition  input  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	410 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	205 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_680_update_completed_
      -- CP-element group 176: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_680_Update/ca
      -- CP-element group 176: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_680_Update/$exit
      -- 
    ca_1389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_680_inst_ack_1, ack => convTranspose_CP_39_elements(176)); -- 
    -- CP-element group 177:  transition  input  output  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	174 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	178 
    -- CP-element group 177:  members (6) 
      -- CP-element group 177: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_689_update_start_
      -- CP-element group 177: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_689_sample_completed_
      -- CP-element group 177: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_689_Update/cr
      -- CP-element group 177: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_689_Update/$entry
      -- CP-element group 177: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_689_Sample/ra
      -- CP-element group 177: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_689_Sample/$exit
      -- 
    ra_1398_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_689_inst_ack_0, ack => convTranspose_CP_39_elements(177)); -- 
    cr_1402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(177), ack => RPIPE_ConvTranspose_input_pipe_689_inst_req_1); -- 
    -- CP-element group 178:  fork  transition  input  output  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	177 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178: 	181 
    -- CP-element group 178:  members (9) 
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_707_Sample/$entry
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_707_Sample/rr
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_707_sample_start_
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_689_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_693_sample_start_
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_689_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_689_Update/ca
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_693_Sample/rr
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_693_Sample/$entry
      -- 
    ca_1403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_689_inst_ack_1, ack => convTranspose_CP_39_elements(178)); -- 
    rr_1425_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1425_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(178), ack => RPIPE_ConvTranspose_input_pipe_707_inst_req_0); -- 
    rr_1411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(178), ack => type_cast_693_inst_req_0); -- 
    -- CP-element group 179:  transition  input  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	178 
    -- CP-element group 179: successors 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_693_sample_completed_
      -- CP-element group 179: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_693_Sample/ra
      -- CP-element group 179: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_693_Sample/$exit
      -- 
    ra_1412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_693_inst_ack_0, ack => convTranspose_CP_39_elements(179)); -- 
    -- CP-element group 180:  transition  input  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	410 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	205 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_693_Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_693_Update/ca
      -- CP-element group 180: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_693_update_completed_
      -- 
    ca_1417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_693_inst_ack_1, ack => convTranspose_CP_39_elements(180)); -- 
    -- CP-element group 181:  transition  input  output  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	178 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	182 
    -- CP-element group 181:  members (6) 
      -- CP-element group 181: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_707_sample_completed_
      -- CP-element group 181: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_707_Sample/$exit
      -- CP-element group 181: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_707_Sample/ra
      -- CP-element group 181: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_707_Update/$entry
      -- CP-element group 181: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_707_update_start_
      -- CP-element group 181: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_707_Update/cr
      -- 
    ra_1426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_707_inst_ack_0, ack => convTranspose_CP_39_elements(181)); -- 
    cr_1430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(181), ack => RPIPE_ConvTranspose_input_pipe_707_inst_req_1); -- 
    -- CP-element group 182:  fork  transition  input  output  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	181 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	185 
    -- CP-element group 182: 	183 
    -- CP-element group 182:  members (9) 
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_711_Sample/rr
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_725_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_725_Sample/rr
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_725_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_711_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_707_update_completed_
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_711_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_707_Update/ca
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_707_Update/$exit
      -- 
    ca_1431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_707_inst_ack_1, ack => convTranspose_CP_39_elements(182)); -- 
    rr_1453_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1453_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(182), ack => RPIPE_ConvTranspose_input_pipe_725_inst_req_0); -- 
    rr_1439_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1439_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(182), ack => type_cast_711_inst_req_0); -- 
    -- CP-element group 183:  transition  input  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	182 
    -- CP-element group 183: successors 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_711_Sample/$exit
      -- CP-element group 183: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_711_Sample/ra
      -- CP-element group 183: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_711_sample_completed_
      -- 
    ra_1440_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_711_inst_ack_0, ack => convTranspose_CP_39_elements(183)); -- 
    -- CP-element group 184:  transition  input  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	410 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	205 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_711_Update/ca
      -- CP-element group 184: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_711_Update/$exit
      -- CP-element group 184: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_711_update_completed_
      -- 
    ca_1445_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_711_inst_ack_1, ack => convTranspose_CP_39_elements(184)); -- 
    -- CP-element group 185:  transition  input  output  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	182 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	186 
    -- CP-element group 185:  members (6) 
      -- CP-element group 185: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_725_Sample/$exit
      -- CP-element group 185: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_725_Sample/ra
      -- CP-element group 185: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_725_update_start_
      -- CP-element group 185: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_725_sample_completed_
      -- CP-element group 185: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_725_Update/$entry
      -- CP-element group 185: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_725_Update/cr
      -- 
    ra_1454_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_725_inst_ack_0, ack => convTranspose_CP_39_elements(185)); -- 
    cr_1458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(185), ack => RPIPE_ConvTranspose_input_pipe_725_inst_req_1); -- 
    -- CP-element group 186:  fork  transition  input  output  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	185 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186: 	189 
    -- CP-element group 186:  members (9) 
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_725_update_completed_
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_725_Update/$exit
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_725_Update/ca
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_729_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_729_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_729_Sample/rr
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_743_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_743_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_743_Sample/rr
      -- 
    ca_1459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_725_inst_ack_1, ack => convTranspose_CP_39_elements(186)); -- 
    rr_1467_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1467_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(186), ack => type_cast_729_inst_req_0); -- 
    rr_1481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(186), ack => RPIPE_ConvTranspose_input_pipe_743_inst_req_0); -- 
    -- CP-element group 187:  transition  input  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_729_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_729_Sample/$exit
      -- CP-element group 187: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_729_Sample/ra
      -- 
    ra_1468_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_729_inst_ack_0, ack => convTranspose_CP_39_elements(187)); -- 
    -- CP-element group 188:  transition  input  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	410 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	205 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_729_update_completed_
      -- CP-element group 188: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_729_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_729_Update/ca
      -- 
    ca_1473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_729_inst_ack_1, ack => convTranspose_CP_39_elements(188)); -- 
    -- CP-element group 189:  transition  input  output  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	186 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	190 
    -- CP-element group 189:  members (6) 
      -- CP-element group 189: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_743_sample_completed_
      -- CP-element group 189: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_743_update_start_
      -- CP-element group 189: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_743_Sample/$exit
      -- CP-element group 189: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_743_Sample/ra
      -- CP-element group 189: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_743_Update/$entry
      -- CP-element group 189: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_743_Update/cr
      -- 
    ra_1482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_743_inst_ack_0, ack => convTranspose_CP_39_elements(189)); -- 
    cr_1486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(189), ack => RPIPE_ConvTranspose_input_pipe_743_inst_req_1); -- 
    -- CP-element group 190:  fork  transition  input  output  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	189 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	191 
    -- CP-element group 190: 	193 
    -- CP-element group 190:  members (9) 
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_743_update_completed_
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_743_Update/$exit
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_743_Update/ca
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_747_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_747_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_747_Sample/rr
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_761_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_761_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_761_Sample/rr
      -- 
    ca_1487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_743_inst_ack_1, ack => convTranspose_CP_39_elements(190)); -- 
    rr_1495_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1495_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(190), ack => type_cast_747_inst_req_0); -- 
    rr_1509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(190), ack => RPIPE_ConvTranspose_input_pipe_761_inst_req_0); -- 
    -- CP-element group 191:  transition  input  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	190 
    -- CP-element group 191: successors 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_747_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_747_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_747_Sample/ra
      -- 
    ra_1496_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_747_inst_ack_0, ack => convTranspose_CP_39_elements(191)); -- 
    -- CP-element group 192:  transition  input  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	410 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	205 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_747_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_747_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_747_Update/ca
      -- 
    ca_1501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_747_inst_ack_1, ack => convTranspose_CP_39_elements(192)); -- 
    -- CP-element group 193:  transition  input  output  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	190 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	194 
    -- CP-element group 193:  members (6) 
      -- CP-element group 193: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_761_sample_completed_
      -- CP-element group 193: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_761_update_start_
      -- CP-element group 193: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_761_Sample/$exit
      -- CP-element group 193: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_761_Sample/ra
      -- CP-element group 193: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_761_Update/$entry
      -- CP-element group 193: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_761_Update/cr
      -- 
    ra_1510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_761_inst_ack_0, ack => convTranspose_CP_39_elements(193)); -- 
    cr_1514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(193), ack => RPIPE_ConvTranspose_input_pipe_761_inst_req_1); -- 
    -- CP-element group 194:  fork  transition  input  output  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	193 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194: 	197 
    -- CP-element group 194:  members (9) 
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_761_update_completed_
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_761_Update/$exit
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_761_Update/ca
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_765_sample_start_
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_765_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_765_Sample/rr
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_779_sample_start_
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_779_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_779_Sample/rr
      -- 
    ca_1515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_761_inst_ack_1, ack => convTranspose_CP_39_elements(194)); -- 
    rr_1523_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1523_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(194), ack => type_cast_765_inst_req_0); -- 
    rr_1537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(194), ack => RPIPE_ConvTranspose_input_pipe_779_inst_req_0); -- 
    -- CP-element group 195:  transition  input  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_765_sample_completed_
      -- CP-element group 195: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_765_Sample/$exit
      -- CP-element group 195: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_765_Sample/ra
      -- 
    ra_1524_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_765_inst_ack_0, ack => convTranspose_CP_39_elements(195)); -- 
    -- CP-element group 196:  transition  input  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	410 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	205 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_765_update_completed_
      -- CP-element group 196: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_765_Update/$exit
      -- CP-element group 196: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_765_Update/ca
      -- 
    ca_1529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_765_inst_ack_1, ack => convTranspose_CP_39_elements(196)); -- 
    -- CP-element group 197:  transition  input  output  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	194 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	198 
    -- CP-element group 197:  members (6) 
      -- CP-element group 197: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_779_sample_completed_
      -- CP-element group 197: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_779_update_start_
      -- CP-element group 197: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_779_Sample/$exit
      -- CP-element group 197: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_779_Sample/ra
      -- CP-element group 197: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_779_Update/$entry
      -- CP-element group 197: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_779_Update/cr
      -- 
    ra_1538_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_779_inst_ack_0, ack => convTranspose_CP_39_elements(197)); -- 
    cr_1542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(197), ack => RPIPE_ConvTranspose_input_pipe_779_inst_req_1); -- 
    -- CP-element group 198:  fork  transition  input  output  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	197 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	199 
    -- CP-element group 198: 	201 
    -- CP-element group 198:  members (9) 
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_779_update_completed_
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_779_Update/$exit
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_779_Update/ca
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_783_sample_start_
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_783_Sample/$entry
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_783_Sample/rr
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_797_sample_start_
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_797_Sample/$entry
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_797_Sample/rr
      -- 
    ca_1543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_779_inst_ack_1, ack => convTranspose_CP_39_elements(198)); -- 
    rr_1551_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1551_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(198), ack => type_cast_783_inst_req_0); -- 
    rr_1565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(198), ack => RPIPE_ConvTranspose_input_pipe_797_inst_req_0); -- 
    -- CP-element group 199:  transition  input  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	198 
    -- CP-element group 199: successors 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_783_sample_completed_
      -- CP-element group 199: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_783_Sample/$exit
      -- CP-element group 199: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_783_Sample/ra
      -- 
    ra_1552_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_783_inst_ack_0, ack => convTranspose_CP_39_elements(199)); -- 
    -- CP-element group 200:  transition  input  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	410 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	205 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_783_update_completed_
      -- CP-element group 200: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_783_Update/$exit
      -- CP-element group 200: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_783_Update/ca
      -- 
    ca_1557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_783_inst_ack_1, ack => convTranspose_CP_39_elements(200)); -- 
    -- CP-element group 201:  transition  input  output  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	198 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201:  members (6) 
      -- CP-element group 201: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_797_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_797_update_start_
      -- CP-element group 201: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_797_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_797_Sample/ra
      -- CP-element group 201: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_797_Update/$entry
      -- CP-element group 201: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_797_Update/cr
      -- 
    ra_1566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_797_inst_ack_0, ack => convTranspose_CP_39_elements(201)); -- 
    cr_1570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(201), ack => RPIPE_ConvTranspose_input_pipe_797_inst_req_1); -- 
    -- CP-element group 202:  transition  input  output  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	201 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202:  members (6) 
      -- CP-element group 202: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_797_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_797_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_797_Update/ca
      -- CP-element group 202: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_801_sample_start_
      -- CP-element group 202: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_801_Sample/$entry
      -- CP-element group 202: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_801_Sample/rr
      -- 
    ca_1571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_797_inst_ack_1, ack => convTranspose_CP_39_elements(202)); -- 
    rr_1579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(202), ack => type_cast_801_inst_req_0); -- 
    -- CP-element group 203:  transition  input  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	202 
    -- CP-element group 203: successors 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_801_sample_completed_
      -- CP-element group 203: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_801_Sample/$exit
      -- CP-element group 203: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_801_Sample/ra
      -- 
    ra_1580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_801_inst_ack_0, ack => convTranspose_CP_39_elements(203)); -- 
    -- CP-element group 204:  transition  input  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	410 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	205 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_801_update_completed_
      -- CP-element group 204: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_801_Update/$exit
      -- CP-element group 204: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_801_Update/ca
      -- 
    ca_1585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_801_inst_ack_1, ack => convTranspose_CP_39_elements(204)); -- 
    -- CP-element group 205:  join  transition  output  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	188 
    -- CP-element group 205: 	192 
    -- CP-element group 205: 	196 
    -- CP-element group 205: 	200 
    -- CP-element group 205: 	204 
    -- CP-element group 205: 	180 
    -- CP-element group 205: 	184 
    -- CP-element group 205: 	172 
    -- CP-element group 205: 	176 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	206 
    -- CP-element group 205:  members (9) 
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_sample_start_
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_Sample/$entry
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_Sample/ptr_deref_809_Split/$entry
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_Sample/ptr_deref_809_Split/$exit
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_Sample/ptr_deref_809_Split/split_req
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_Sample/ptr_deref_809_Split/split_ack
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_Sample/word_access_start/$entry
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_Sample/word_access_start/word_0/$entry
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_Sample/word_access_start/word_0/rr
      -- 
    rr_1623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(205), ack => ptr_deref_809_store_0_req_0); -- 
    convTranspose_cp_element_group_205: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_205"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(188) & convTranspose_CP_39_elements(192) & convTranspose_CP_39_elements(196) & convTranspose_CP_39_elements(200) & convTranspose_CP_39_elements(204) & convTranspose_CP_39_elements(180) & convTranspose_CP_39_elements(184) & convTranspose_CP_39_elements(172) & convTranspose_CP_39_elements(176);
      gj_convTranspose_cp_element_group_205 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(205), clk => clk, reset => reset); --
    end block;
    -- CP-element group 206:  transition  input  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	205 
    -- CP-element group 206: successors 
    -- CP-element group 206:  members (5) 
      -- CP-element group 206: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_sample_completed_
      -- CP-element group 206: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_Sample/$exit
      -- CP-element group 206: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_Sample/word_access_start/$exit
      -- CP-element group 206: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_Sample/word_access_start/word_0/$exit
      -- CP-element group 206: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_Sample/word_access_start/word_0/ra
      -- 
    ra_1624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_809_store_0_ack_0, ack => convTranspose_CP_39_elements(206)); -- 
    -- CP-element group 207:  transition  input  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	410 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	208 
    -- CP-element group 207:  members (5) 
      -- CP-element group 207: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_update_completed_
      -- CP-element group 207: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_Update/$exit
      -- CP-element group 207: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_Update/word_access_complete/$exit
      -- CP-element group 207: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_Update/word_access_complete/word_0/$exit
      -- CP-element group 207: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_Update/word_access_complete/word_0/ca
      -- 
    ca_1635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_809_store_0_ack_1, ack => convTranspose_CP_39_elements(207)); -- 
    -- CP-element group 208:  branch  join  transition  place  output  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	207 
    -- CP-element group 208: 	169 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	209 
    -- CP-element group 208: 	210 
    -- CP-element group 208:  members (10) 
      -- CP-element group 208: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822__exit__
      -- CP-element group 208: 	 branch_block_stmt_33/if_stmt_823__entry__
      -- CP-element group 208: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/$exit
      -- CP-element group 208: 	 branch_block_stmt_33/if_stmt_823_dead_link/$entry
      -- CP-element group 208: 	 branch_block_stmt_33/if_stmt_823_eval_test/$entry
      -- CP-element group 208: 	 branch_block_stmt_33/if_stmt_823_eval_test/$exit
      -- CP-element group 208: 	 branch_block_stmt_33/if_stmt_823_eval_test/branch_req
      -- CP-element group 208: 	 branch_block_stmt_33/R_exitcond2_824_place
      -- CP-element group 208: 	 branch_block_stmt_33/if_stmt_823_if_link/$entry
      -- CP-element group 208: 	 branch_block_stmt_33/if_stmt_823_else_link/$entry
      -- 
    branch_req_1643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(208), ack => if_stmt_823_branch_req_0); -- 
    convTranspose_cp_element_group_208: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_208"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(207) & convTranspose_CP_39_elements(169);
      gj_convTranspose_cp_element_group_208 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(208), clk => clk, reset => reset); --
    end block;
    -- CP-element group 209:  merge  transition  place  input  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	208 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	411 
    -- CP-element group 209:  members (13) 
      -- CP-element group 209: 	 branch_block_stmt_33/merge_stmt_829__exit__
      -- CP-element group 209: 	 branch_block_stmt_33/forx_xend236x_xloopexit_forx_xend236
      -- CP-element group 209: 	 branch_block_stmt_33/merge_stmt_829_PhiReqMerge
      -- CP-element group 209: 	 branch_block_stmt_33/if_stmt_823_if_link/$exit
      -- CP-element group 209: 	 branch_block_stmt_33/if_stmt_823_if_link/if_choice_transition
      -- CP-element group 209: 	 branch_block_stmt_33/forx_xbody182_forx_xend236x_xloopexit
      -- CP-element group 209: 	 branch_block_stmt_33/forx_xend236x_xloopexit_forx_xend236_PhiReq/$exit
      -- CP-element group 209: 	 branch_block_stmt_33/forx_xend236x_xloopexit_forx_xend236_PhiReq/$entry
      -- CP-element group 209: 	 branch_block_stmt_33/merge_stmt_829_PhiAck/dummy
      -- CP-element group 209: 	 branch_block_stmt_33/merge_stmt_829_PhiAck/$exit
      -- CP-element group 209: 	 branch_block_stmt_33/merge_stmt_829_PhiAck/$entry
      -- CP-element group 209: 	 branch_block_stmt_33/forx_xbody182_forx_xend236x_xloopexit_PhiReq/$exit
      -- CP-element group 209: 	 branch_block_stmt_33/forx_xbody182_forx_xend236x_xloopexit_PhiReq/$entry
      -- 
    if_choice_transition_1648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_823_branch_ack_1, ack => convTranspose_CP_39_elements(209)); -- 
    -- CP-element group 210:  fork  transition  place  input  output  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	208 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	406 
    -- CP-element group 210: 	407 
    -- CP-element group 210:  members (12) 
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_660/phi_stmt_660_sources/type_cast_663/SplitProtocol/Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_33/if_stmt_823_else_link/$exit
      -- CP-element group 210: 	 branch_block_stmt_33/if_stmt_823_else_link/else_choice_transition
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody182_forx_xbody182
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_660/phi_stmt_660_sources/type_cast_663/SplitProtocol/$entry
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_660/phi_stmt_660_sources/type_cast_663/SplitProtocol/Sample/rr
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_660/phi_stmt_660_sources/type_cast_663/SplitProtocol/Update/$entry
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_660/phi_stmt_660_sources/type_cast_663/SplitProtocol/Update/cr
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody182_forx_xbody182_PhiReq/$entry
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_660/phi_stmt_660_sources/type_cast_663/$entry
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_660/phi_stmt_660_sources/$entry
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_660/$entry
      -- 
    else_choice_transition_1652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_823_branch_ack_0, ack => convTranspose_CP_39_elements(210)); -- 
    rr_3154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(210), ack => type_cast_663_inst_req_0); -- 
    cr_3159_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3159_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(210), ack => type_cast_663_inst_req_1); -- 
    -- CP-element group 211:  transition  input  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	411 
    -- CP-element group 211: successors 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_834_sample_completed_
      -- CP-element group 211: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_834_Sample/$exit
      -- CP-element group 211: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_834_Sample/ra
      -- 
    ra_1666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_834_inst_ack_0, ack => convTranspose_CP_39_elements(211)); -- 
    -- CP-element group 212:  transition  input  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	411 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	217 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_834_update_completed_
      -- CP-element group 212: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_834_Update/$exit
      -- CP-element group 212: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_834_Update/ca
      -- 
    ca_1671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_834_inst_ack_1, ack => convTranspose_CP_39_elements(212)); -- 
    -- CP-element group 213:  transition  input  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	411 
    -- CP-element group 213: successors 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_838_sample_completed_
      -- CP-element group 213: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_838_Sample/$exit
      -- CP-element group 213: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_838_Sample/ra
      -- 
    ra_1680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_838_inst_ack_0, ack => convTranspose_CP_39_elements(213)); -- 
    -- CP-element group 214:  transition  input  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	411 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	217 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_838_update_completed_
      -- CP-element group 214: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_838_Update/$exit
      -- CP-element group 214: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_838_Update/ca
      -- 
    ca_1685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_838_inst_ack_1, ack => convTranspose_CP_39_elements(214)); -- 
    -- CP-element group 215:  transition  input  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	411 
    -- CP-element group 215: successors 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_842_sample_completed_
      -- CP-element group 215: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_842_Sample/$exit
      -- CP-element group 215: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_842_Sample/ra
      -- 
    ra_1694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_842_inst_ack_0, ack => convTranspose_CP_39_elements(215)); -- 
    -- CP-element group 216:  transition  input  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	411 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	217 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_842_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_842_Update/$exit
      -- CP-element group 216: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_842_Update/ca
      -- 
    ca_1699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_842_inst_ack_1, ack => convTranspose_CP_39_elements(216)); -- 
    -- CP-element group 217:  branch  join  transition  place  output  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	212 
    -- CP-element group 217: 	214 
    -- CP-element group 217: 	216 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	218 
    -- CP-element group 217: 	219 
    -- CP-element group 217:  members (10) 
      -- CP-element group 217: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859__exit__
      -- CP-element group 217: 	 branch_block_stmt_33/if_stmt_860__entry__
      -- CP-element group 217: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/$exit
      -- CP-element group 217: 	 branch_block_stmt_33/if_stmt_860_dead_link/$entry
      -- CP-element group 217: 	 branch_block_stmt_33/if_stmt_860_eval_test/$entry
      -- CP-element group 217: 	 branch_block_stmt_33/if_stmt_860_eval_test/$exit
      -- CP-element group 217: 	 branch_block_stmt_33/if_stmt_860_eval_test/branch_req
      -- CP-element group 217: 	 branch_block_stmt_33/R_cmp250409_861_place
      -- CP-element group 217: 	 branch_block_stmt_33/if_stmt_860_if_link/$entry
      -- CP-element group 217: 	 branch_block_stmt_33/if_stmt_860_else_link/$entry
      -- 
    branch_req_1707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(217), ack => if_stmt_860_branch_req_0); -- 
    convTranspose_cp_element_group_217: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_217"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(212) & convTranspose_CP_39_elements(214) & convTranspose_CP_39_elements(216);
      gj_convTranspose_cp_element_group_217 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(217), clk => clk, reset => reset); --
    end block;
    -- CP-element group 218:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	217 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	220 
    -- CP-element group 218: 	221 
    -- CP-element group 218:  members (18) 
      -- CP-element group 218: 	 branch_block_stmt_33/merge_stmt_866__exit__
      -- CP-element group 218: 	 branch_block_stmt_33/assign_stmt_872_to_assign_stmt_901__entry__
      -- CP-element group 218: 	 branch_block_stmt_33/merge_stmt_866_PhiReqMerge
      -- CP-element group 218: 	 branch_block_stmt_33/if_stmt_860_if_link/$exit
      -- CP-element group 218: 	 branch_block_stmt_33/if_stmt_860_if_link/if_choice_transition
      -- CP-element group 218: 	 branch_block_stmt_33/forx_xend236_bbx_xnph411
      -- CP-element group 218: 	 branch_block_stmt_33/assign_stmt_872_to_assign_stmt_901/$entry
      -- CP-element group 218: 	 branch_block_stmt_33/assign_stmt_872_to_assign_stmt_901/type_cast_887_sample_start_
      -- CP-element group 218: 	 branch_block_stmt_33/assign_stmt_872_to_assign_stmt_901/type_cast_887_update_start_
      -- CP-element group 218: 	 branch_block_stmt_33/assign_stmt_872_to_assign_stmt_901/type_cast_887_Sample/$entry
      -- CP-element group 218: 	 branch_block_stmt_33/assign_stmt_872_to_assign_stmt_901/type_cast_887_Sample/rr
      -- CP-element group 218: 	 branch_block_stmt_33/assign_stmt_872_to_assign_stmt_901/type_cast_887_Update/$entry
      -- CP-element group 218: 	 branch_block_stmt_33/assign_stmt_872_to_assign_stmt_901/type_cast_887_Update/cr
      -- CP-element group 218: 	 branch_block_stmt_33/merge_stmt_866_PhiAck/dummy
      -- CP-element group 218: 	 branch_block_stmt_33/merge_stmt_866_PhiAck/$exit
      -- CP-element group 218: 	 branch_block_stmt_33/merge_stmt_866_PhiAck/$entry
      -- CP-element group 218: 	 branch_block_stmt_33/forx_xend236_bbx_xnph411_PhiReq/$exit
      -- CP-element group 218: 	 branch_block_stmt_33/forx_xend236_bbx_xnph411_PhiReq/$entry
      -- 
    if_choice_transition_1712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_860_branch_ack_1, ack => convTranspose_CP_39_elements(218)); -- 
    rr_1729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(218), ack => type_cast_887_inst_req_0); -- 
    cr_1734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(218), ack => type_cast_887_inst_req_1); -- 
    -- CP-element group 219:  transition  place  input  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	217 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	418 
    -- CP-element group 219:  members (5) 
      -- CP-element group 219: 	 branch_block_stmt_33/if_stmt_860_else_link/$exit
      -- CP-element group 219: 	 branch_block_stmt_33/if_stmt_860_else_link/else_choice_transition
      -- CP-element group 219: 	 branch_block_stmt_33/forx_xend236_forx_xend259
      -- CP-element group 219: 	 branch_block_stmt_33/forx_xend236_forx_xend259_PhiReq/$exit
      -- CP-element group 219: 	 branch_block_stmt_33/forx_xend236_forx_xend259_PhiReq/$entry
      -- 
    else_choice_transition_1716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_860_branch_ack_0, ack => convTranspose_CP_39_elements(219)); -- 
    -- CP-element group 220:  transition  input  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	218 
    -- CP-element group 220: successors 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_33/assign_stmt_872_to_assign_stmt_901/type_cast_887_sample_completed_
      -- CP-element group 220: 	 branch_block_stmt_33/assign_stmt_872_to_assign_stmt_901/type_cast_887_Sample/$exit
      -- CP-element group 220: 	 branch_block_stmt_33/assign_stmt_872_to_assign_stmt_901/type_cast_887_Sample/ra
      -- 
    ra_1730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_887_inst_ack_0, ack => convTranspose_CP_39_elements(220)); -- 
    -- CP-element group 221:  transition  place  input  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	218 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	412 
    -- CP-element group 221:  members (9) 
      -- CP-element group 221: 	 branch_block_stmt_33/assign_stmt_872_to_assign_stmt_901__exit__
      -- CP-element group 221: 	 branch_block_stmt_33/bbx_xnph411_forx_xbody252
      -- CP-element group 221: 	 branch_block_stmt_33/assign_stmt_872_to_assign_stmt_901/$exit
      -- CP-element group 221: 	 branch_block_stmt_33/assign_stmt_872_to_assign_stmt_901/type_cast_887_update_completed_
      -- CP-element group 221: 	 branch_block_stmt_33/assign_stmt_872_to_assign_stmt_901/type_cast_887_Update/$exit
      -- CP-element group 221: 	 branch_block_stmt_33/assign_stmt_872_to_assign_stmt_901/type_cast_887_Update/ca
      -- CP-element group 221: 	 branch_block_stmt_33/bbx_xnph411_forx_xbody252_PhiReq/phi_stmt_904/phi_stmt_904_sources/$entry
      -- CP-element group 221: 	 branch_block_stmt_33/bbx_xnph411_forx_xbody252_PhiReq/phi_stmt_904/$entry
      -- CP-element group 221: 	 branch_block_stmt_33/bbx_xnph411_forx_xbody252_PhiReq/$entry
      -- 
    ca_1735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_887_inst_ack_1, ack => convTranspose_CP_39_elements(221)); -- 
    -- CP-element group 222:  transition  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	417 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	228 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_final_index_sum_regn_sample_complete
      -- CP-element group 222: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_final_index_sum_regn_Sample/$exit
      -- CP-element group 222: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_final_index_sum_regn_Sample/ack
      -- 
    ack_1764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_916_index_offset_ack_0, ack => convTranspose_CP_39_elements(222)); -- 
    -- CP-element group 223:  transition  input  output  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	417 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223:  members (11) 
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/addr_of_917_sample_start_
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_root_address_calculated
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_offset_calculated
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_final_index_sum_regn_Update/$exit
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_final_index_sum_regn_Update/ack
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_base_plus_offset/$entry
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_base_plus_offset/$exit
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_base_plus_offset/sum_rename_req
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_base_plus_offset/sum_rename_ack
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/addr_of_917_request/$entry
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/addr_of_917_request/req
      -- 
    ack_1769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_916_index_offset_ack_1, ack => convTranspose_CP_39_elements(223)); -- 
    req_1778_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1778_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(223), ack => addr_of_917_final_reg_req_0); -- 
    -- CP-element group 224:  transition  input  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/addr_of_917_sample_completed_
      -- CP-element group 224: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/addr_of_917_request/$exit
      -- CP-element group 224: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/addr_of_917_request/ack
      -- 
    ack_1779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_917_final_reg_ack_0, ack => convTranspose_CP_39_elements(224)); -- 
    -- CP-element group 225:  join  fork  transition  input  output  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	417 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	226 
    -- CP-element group 225:  members (28) 
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/addr_of_917_update_completed_
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/addr_of_917_complete/$exit
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/addr_of_917_complete/ack
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_sample_start_
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_base_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_word_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_root_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_base_address_resized
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_base_addr_resize/$entry
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_base_addr_resize/$exit
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_base_addr_resize/base_resize_req
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_base_addr_resize/base_resize_ack
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_base_plus_offset/$entry
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_base_plus_offset/$exit
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_base_plus_offset/sum_rename_req
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_base_plus_offset/sum_rename_ack
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_word_addrgen/$entry
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_word_addrgen/$exit
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_word_addrgen/root_register_req
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_word_addrgen/root_register_ack
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_Sample/$entry
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_Sample/ptr_deref_920_Split/$entry
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_Sample/ptr_deref_920_Split/$exit
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_Sample/ptr_deref_920_Split/split_req
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_Sample/ptr_deref_920_Split/split_ack
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_Sample/word_access_start/$entry
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_Sample/word_access_start/word_0/$entry
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_Sample/word_access_start/word_0/rr
      -- 
    ack_1784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_917_final_reg_ack_1, ack => convTranspose_CP_39_elements(225)); -- 
    rr_1822_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1822_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(225), ack => ptr_deref_920_store_0_req_0); -- 
    -- CP-element group 226:  transition  input  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	225 
    -- CP-element group 226: successors 
    -- CP-element group 226:  members (5) 
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_sample_completed_
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_Sample/$exit
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_Sample/word_access_start/$exit
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_Sample/word_access_start/word_0/$exit
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_Sample/word_access_start/word_0/ra
      -- 
    ra_1823_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_920_store_0_ack_0, ack => convTranspose_CP_39_elements(226)); -- 
    -- CP-element group 227:  transition  input  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	417 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	228 
    -- CP-element group 227:  members (5) 
      -- CP-element group 227: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_update_completed_
      -- CP-element group 227: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_Update/$exit
      -- CP-element group 227: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_Update/word_access_complete/$exit
      -- CP-element group 227: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_Update/word_access_complete/word_0/$exit
      -- CP-element group 227: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_Update/word_access_complete/word_0/ca
      -- 
    ca_1834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_920_store_0_ack_1, ack => convTranspose_CP_39_elements(227)); -- 
    -- CP-element group 228:  branch  join  transition  place  output  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	222 
    -- CP-element group 228: 	227 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	229 
    -- CP-element group 228: 	230 
    -- CP-element group 228:  members (10) 
      -- CP-element group 228: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934__exit__
      -- CP-element group 228: 	 branch_block_stmt_33/if_stmt_935__entry__
      -- CP-element group 228: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/$exit
      -- CP-element group 228: 	 branch_block_stmt_33/if_stmt_935_dead_link/$entry
      -- CP-element group 228: 	 branch_block_stmt_33/if_stmt_935_eval_test/$entry
      -- CP-element group 228: 	 branch_block_stmt_33/if_stmt_935_eval_test/$exit
      -- CP-element group 228: 	 branch_block_stmt_33/if_stmt_935_eval_test/branch_req
      -- CP-element group 228: 	 branch_block_stmt_33/R_exitcond_936_place
      -- CP-element group 228: 	 branch_block_stmt_33/if_stmt_935_if_link/$entry
      -- CP-element group 228: 	 branch_block_stmt_33/if_stmt_935_else_link/$entry
      -- 
    branch_req_1842_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1842_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(228), ack => if_stmt_935_branch_req_0); -- 
    convTranspose_cp_element_group_228: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_228"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(222) & convTranspose_CP_39_elements(227);
      gj_convTranspose_cp_element_group_228 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(228), clk => clk, reset => reset); --
    end block;
    -- CP-element group 229:  merge  transition  place  input  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	228 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	418 
    -- CP-element group 229:  members (13) 
      -- CP-element group 229: 	 branch_block_stmt_33/merge_stmt_941__exit__
      -- CP-element group 229: 	 branch_block_stmt_33/forx_xend259x_xloopexit_forx_xend259
      -- CP-element group 229: 	 branch_block_stmt_33/merge_stmt_941_PhiReqMerge
      -- CP-element group 229: 	 branch_block_stmt_33/if_stmt_935_if_link/$exit
      -- CP-element group 229: 	 branch_block_stmt_33/if_stmt_935_if_link/if_choice_transition
      -- CP-element group 229: 	 branch_block_stmt_33/forx_xbody252_forx_xend259x_xloopexit
      -- CP-element group 229: 	 branch_block_stmt_33/forx_xend259x_xloopexit_forx_xend259_PhiReq/$exit
      -- CP-element group 229: 	 branch_block_stmt_33/forx_xend259x_xloopexit_forx_xend259_PhiReq/$entry
      -- CP-element group 229: 	 branch_block_stmt_33/merge_stmt_941_PhiAck/dummy
      -- CP-element group 229: 	 branch_block_stmt_33/merge_stmt_941_PhiAck/$exit
      -- CP-element group 229: 	 branch_block_stmt_33/merge_stmt_941_PhiAck/$entry
      -- CP-element group 229: 	 branch_block_stmt_33/forx_xbody252_forx_xend259x_xloopexit_PhiReq/$exit
      -- CP-element group 229: 	 branch_block_stmt_33/forx_xbody252_forx_xend259x_xloopexit_PhiReq/$entry
      -- 
    if_choice_transition_1847_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_935_branch_ack_1, ack => convTranspose_CP_39_elements(229)); -- 
    -- CP-element group 230:  fork  transition  place  input  output  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	228 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	413 
    -- CP-element group 230: 	414 
    -- CP-element group 230:  members (12) 
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody252_forx_xbody252_PhiReq/phi_stmt_904/phi_stmt_904_sources/type_cast_910/SplitProtocol/$entry
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody252_forx_xbody252_PhiReq/phi_stmt_904/phi_stmt_904_sources/type_cast_910/SplitProtocol/Sample/rr
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody252_forx_xbody252_PhiReq/phi_stmt_904/phi_stmt_904_sources/type_cast_910/SplitProtocol/Sample/$entry
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody252_forx_xbody252_PhiReq/phi_stmt_904/phi_stmt_904_sources/type_cast_910/$entry
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody252_forx_xbody252_PhiReq/phi_stmt_904/phi_stmt_904_sources/$entry
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody252_forx_xbody252_PhiReq/phi_stmt_904/phi_stmt_904_sources/type_cast_910/SplitProtocol/Update/$entry
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody252_forx_xbody252_PhiReq/phi_stmt_904/phi_stmt_904_sources/type_cast_910/SplitProtocol/Update/cr
      -- CP-element group 230: 	 branch_block_stmt_33/if_stmt_935_else_link/$exit
      -- CP-element group 230: 	 branch_block_stmt_33/if_stmt_935_else_link/else_choice_transition
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody252_forx_xbody252
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody252_forx_xbody252_PhiReq/phi_stmt_904/$entry
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody252_forx_xbody252_PhiReq/$entry
      -- 
    else_choice_transition_1851_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_935_branch_ack_0, ack => convTranspose_CP_39_elements(230)); -- 
    rr_3231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(230), ack => type_cast_910_inst_req_0); -- 
    cr_3236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(230), ack => type_cast_910_inst_req_1); -- 
    -- CP-element group 231:  transition  input  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	418 
    -- CP-element group 231: successors 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/call_stmt_946_sample_completed_
      -- CP-element group 231: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/call_stmt_946_Sample/$exit
      -- CP-element group 231: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/call_stmt_946_Sample/cra
      -- 
    cra_1865_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_946_call_ack_0, ack => convTranspose_CP_39_elements(231)); -- 
    -- CP-element group 232:  transition  input  output  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	418 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	233 
    -- CP-element group 232:  members (6) 
      -- CP-element group 232: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/call_stmt_946_update_completed_
      -- CP-element group 232: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/call_stmt_946_Update/$exit
      -- CP-element group 232: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/call_stmt_946_Update/cca
      -- CP-element group 232: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/type_cast_951_sample_start_
      -- CP-element group 232: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/type_cast_951_Sample/$entry
      -- CP-element group 232: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/type_cast_951_Sample/rr
      -- 
    cca_1870_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_946_call_ack_1, ack => convTranspose_CP_39_elements(232)); -- 
    rr_1878_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1878_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(232), ack => type_cast_951_inst_req_0); -- 
    -- CP-element group 233:  transition  input  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	232 
    -- CP-element group 233: successors 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/type_cast_951_sample_completed_
      -- CP-element group 233: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/type_cast_951_Sample/$exit
      -- CP-element group 233: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/type_cast_951_Sample/ra
      -- 
    ra_1879_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_951_inst_ack_0, ack => convTranspose_CP_39_elements(233)); -- 
    -- CP-element group 234:  transition  input  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	418 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	339 
    -- CP-element group 234:  members (3) 
      -- CP-element group 234: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/type_cast_951_update_completed_
      -- CP-element group 234: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/type_cast_951_Update/$exit
      -- CP-element group 234: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/type_cast_951_Update/ca
      -- 
    ca_1884_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_951_inst_ack_1, ack => convTranspose_CP_39_elements(234)); -- 
    -- CP-element group 235:  transition  input  output  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	418 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235:  members (6) 
      -- CP-element group 235: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_953_sample_completed_
      -- CP-element group 235: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_953_update_start_
      -- CP-element group 235: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_953_Sample/$exit
      -- CP-element group 235: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_953_Sample/ack
      -- CP-element group 235: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_953_Update/$entry
      -- CP-element group 235: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_953_Update/req
      -- 
    ack_1893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_953_inst_ack_0, ack => convTranspose_CP_39_elements(235)); -- 
    req_1897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(235), ack => WPIPE_Block0_start_953_inst_req_1); -- 
    -- CP-element group 236:  transition  input  output  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	237 
    -- CP-element group 236:  members (6) 
      -- CP-element group 236: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_953_update_completed_
      -- CP-element group 236: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_953_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_953_Update/ack
      -- CP-element group 236: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_956_sample_start_
      -- CP-element group 236: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_956_Sample/$entry
      -- CP-element group 236: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_956_Sample/req
      -- 
    ack_1898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_953_inst_ack_1, ack => convTranspose_CP_39_elements(236)); -- 
    req_1906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(236), ack => WPIPE_Block0_start_956_inst_req_0); -- 
    -- CP-element group 237:  transition  input  output  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	236 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	238 
    -- CP-element group 237:  members (6) 
      -- CP-element group 237: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_956_sample_completed_
      -- CP-element group 237: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_956_update_start_
      -- CP-element group 237: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_956_Sample/$exit
      -- CP-element group 237: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_956_Sample/ack
      -- CP-element group 237: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_956_Update/$entry
      -- CP-element group 237: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_956_Update/req
      -- 
    ack_1907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_956_inst_ack_0, ack => convTranspose_CP_39_elements(237)); -- 
    req_1911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(237), ack => WPIPE_Block0_start_956_inst_req_1); -- 
    -- CP-element group 238:  transition  input  output  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	237 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	239 
    -- CP-element group 238:  members (6) 
      -- CP-element group 238: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_956_update_completed_
      -- CP-element group 238: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_956_Update/$exit
      -- CP-element group 238: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_956_Update/ack
      -- CP-element group 238: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_959_sample_start_
      -- CP-element group 238: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_959_Sample/$entry
      -- CP-element group 238: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_959_Sample/req
      -- 
    ack_1912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_956_inst_ack_1, ack => convTranspose_CP_39_elements(238)); -- 
    req_1920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(238), ack => WPIPE_Block0_start_959_inst_req_0); -- 
    -- CP-element group 239:  transition  input  output  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	238 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	240 
    -- CP-element group 239:  members (6) 
      -- CP-element group 239: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_959_sample_completed_
      -- CP-element group 239: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_959_update_start_
      -- CP-element group 239: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_959_Sample/$exit
      -- CP-element group 239: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_959_Sample/ack
      -- CP-element group 239: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_959_Update/$entry
      -- CP-element group 239: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_959_Update/req
      -- 
    ack_1921_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_959_inst_ack_0, ack => convTranspose_CP_39_elements(239)); -- 
    req_1925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(239), ack => WPIPE_Block0_start_959_inst_req_1); -- 
    -- CP-element group 240:  transition  input  output  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	239 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	241 
    -- CP-element group 240:  members (6) 
      -- CP-element group 240: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_959_update_completed_
      -- CP-element group 240: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_959_Update/$exit
      -- CP-element group 240: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_959_Update/ack
      -- CP-element group 240: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_962_sample_start_
      -- CP-element group 240: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_962_Sample/$entry
      -- CP-element group 240: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_962_Sample/req
      -- 
    ack_1926_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_959_inst_ack_1, ack => convTranspose_CP_39_elements(240)); -- 
    req_1934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(240), ack => WPIPE_Block0_start_962_inst_req_0); -- 
    -- CP-element group 241:  transition  input  output  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	240 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	242 
    -- CP-element group 241:  members (6) 
      -- CP-element group 241: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_962_sample_completed_
      -- CP-element group 241: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_962_update_start_
      -- CP-element group 241: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_962_Sample/$exit
      -- CP-element group 241: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_962_Sample/ack
      -- CP-element group 241: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_962_Update/$entry
      -- CP-element group 241: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_962_Update/req
      -- 
    ack_1935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_962_inst_ack_0, ack => convTranspose_CP_39_elements(241)); -- 
    req_1939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(241), ack => WPIPE_Block0_start_962_inst_req_1); -- 
    -- CP-element group 242:  transition  input  output  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	241 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	243 
    -- CP-element group 242:  members (6) 
      -- CP-element group 242: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_962_update_completed_
      -- CP-element group 242: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_962_Update/$exit
      -- CP-element group 242: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_962_Update/ack
      -- CP-element group 242: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_965_sample_start_
      -- CP-element group 242: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_965_Sample/$entry
      -- CP-element group 242: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_965_Sample/req
      -- 
    ack_1940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_962_inst_ack_1, ack => convTranspose_CP_39_elements(242)); -- 
    req_1948_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1948_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(242), ack => WPIPE_Block0_start_965_inst_req_0); -- 
    -- CP-element group 243:  transition  input  output  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	242 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	244 
    -- CP-element group 243:  members (6) 
      -- CP-element group 243: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_965_sample_completed_
      -- CP-element group 243: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_965_update_start_
      -- CP-element group 243: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_965_Sample/$exit
      -- CP-element group 243: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_965_Sample/ack
      -- CP-element group 243: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_965_Update/$entry
      -- CP-element group 243: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_965_Update/req
      -- 
    ack_1949_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_965_inst_ack_0, ack => convTranspose_CP_39_elements(243)); -- 
    req_1953_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1953_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(243), ack => WPIPE_Block0_start_965_inst_req_1); -- 
    -- CP-element group 244:  transition  input  output  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	243 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	245 
    -- CP-element group 244:  members (6) 
      -- CP-element group 244: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_965_update_completed_
      -- CP-element group 244: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_965_Update/$exit
      -- CP-element group 244: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_965_Update/ack
      -- CP-element group 244: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_968_sample_start_
      -- CP-element group 244: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_968_Sample/$entry
      -- CP-element group 244: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_968_Sample/req
      -- 
    ack_1954_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_965_inst_ack_1, ack => convTranspose_CP_39_elements(244)); -- 
    req_1962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(244), ack => WPIPE_Block0_start_968_inst_req_0); -- 
    -- CP-element group 245:  transition  input  output  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	244 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	246 
    -- CP-element group 245:  members (6) 
      -- CP-element group 245: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_968_sample_completed_
      -- CP-element group 245: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_968_update_start_
      -- CP-element group 245: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_968_Sample/$exit
      -- CP-element group 245: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_968_Sample/ack
      -- CP-element group 245: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_968_Update/$entry
      -- CP-element group 245: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_968_Update/req
      -- 
    ack_1963_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_968_inst_ack_0, ack => convTranspose_CP_39_elements(245)); -- 
    req_1967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(245), ack => WPIPE_Block0_start_968_inst_req_1); -- 
    -- CP-element group 246:  transition  input  output  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	245 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	247 
    -- CP-element group 246:  members (6) 
      -- CP-element group 246: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_968_update_completed_
      -- CP-element group 246: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_968_Update/$exit
      -- CP-element group 246: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_968_Update/ack
      -- CP-element group 246: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_971_sample_start_
      -- CP-element group 246: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_971_Sample/$entry
      -- CP-element group 246: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_971_Sample/req
      -- 
    ack_1968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_968_inst_ack_1, ack => convTranspose_CP_39_elements(246)); -- 
    req_1976_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1976_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(246), ack => WPIPE_Block0_start_971_inst_req_0); -- 
    -- CP-element group 247:  transition  input  output  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	246 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	248 
    -- CP-element group 247:  members (6) 
      -- CP-element group 247: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_971_sample_completed_
      -- CP-element group 247: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_971_update_start_
      -- CP-element group 247: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_971_Sample/$exit
      -- CP-element group 247: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_971_Sample/ack
      -- CP-element group 247: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_971_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_971_Update/req
      -- 
    ack_1977_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_971_inst_ack_0, ack => convTranspose_CP_39_elements(247)); -- 
    req_1981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(247), ack => WPIPE_Block0_start_971_inst_req_1); -- 
    -- CP-element group 248:  transition  input  output  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	247 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	249 
    -- CP-element group 248:  members (6) 
      -- CP-element group 248: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_971_update_completed_
      -- CP-element group 248: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_971_Update/$exit
      -- CP-element group 248: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_971_Update/ack
      -- CP-element group 248: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_974_sample_start_
      -- CP-element group 248: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_974_Sample/$entry
      -- CP-element group 248: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_974_Sample/req
      -- 
    ack_1982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_971_inst_ack_1, ack => convTranspose_CP_39_elements(248)); -- 
    req_1990_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1990_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(248), ack => WPIPE_Block0_start_974_inst_req_0); -- 
    -- CP-element group 249:  transition  input  output  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	248 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	250 
    -- CP-element group 249:  members (6) 
      -- CP-element group 249: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_974_sample_completed_
      -- CP-element group 249: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_974_update_start_
      -- CP-element group 249: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_974_Sample/$exit
      -- CP-element group 249: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_974_Sample/ack
      -- CP-element group 249: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_974_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_974_Update/req
      -- 
    ack_1991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_974_inst_ack_0, ack => convTranspose_CP_39_elements(249)); -- 
    req_1995_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1995_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(249), ack => WPIPE_Block0_start_974_inst_req_1); -- 
    -- CP-element group 250:  transition  input  output  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	249 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	251 
    -- CP-element group 250:  members (6) 
      -- CP-element group 250: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_974_update_completed_
      -- CP-element group 250: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_974_Update/$exit
      -- CP-element group 250: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_974_Update/ack
      -- CP-element group 250: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_977_sample_start_
      -- CP-element group 250: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_977_Sample/$entry
      -- CP-element group 250: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_977_Sample/req
      -- 
    ack_1996_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_974_inst_ack_1, ack => convTranspose_CP_39_elements(250)); -- 
    req_2004_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2004_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(250), ack => WPIPE_Block0_start_977_inst_req_0); -- 
    -- CP-element group 251:  transition  input  output  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	250 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	252 
    -- CP-element group 251:  members (6) 
      -- CP-element group 251: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_977_Update/req
      -- CP-element group 251: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_977_Update/$entry
      -- CP-element group 251: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_977_sample_completed_
      -- CP-element group 251: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_977_update_start_
      -- CP-element group 251: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_977_Sample/$exit
      -- CP-element group 251: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_977_Sample/ack
      -- 
    ack_2005_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_977_inst_ack_0, ack => convTranspose_CP_39_elements(251)); -- 
    req_2009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(251), ack => WPIPE_Block0_start_977_inst_req_1); -- 
    -- CP-element group 252:  transition  input  output  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	251 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	253 
    -- CP-element group 252:  members (6) 
      -- CP-element group 252: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_980_Sample/req
      -- CP-element group 252: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_980_Sample/$entry
      -- CP-element group 252: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_980_sample_start_
      -- CP-element group 252: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_977_Update/ack
      -- CP-element group 252: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_977_Update/$exit
      -- CP-element group 252: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_977_update_completed_
      -- 
    ack_2010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_977_inst_ack_1, ack => convTranspose_CP_39_elements(252)); -- 
    req_2018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(252), ack => WPIPE_Block0_start_980_inst_req_0); -- 
    -- CP-element group 253:  transition  input  output  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	252 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	254 
    -- CP-element group 253:  members (6) 
      -- CP-element group 253: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_980_update_start_
      -- CP-element group 253: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_980_sample_completed_
      -- CP-element group 253: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_980_Sample/ack
      -- CP-element group 253: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_980_Update/$entry
      -- CP-element group 253: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_980_Update/req
      -- CP-element group 253: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_980_Sample/$exit
      -- 
    ack_2019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_980_inst_ack_0, ack => convTranspose_CP_39_elements(253)); -- 
    req_2023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(253), ack => WPIPE_Block0_start_980_inst_req_1); -- 
    -- CP-element group 254:  transition  input  output  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	253 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	255 
    -- CP-element group 254:  members (6) 
      -- CP-element group 254: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_980_update_completed_
      -- CP-element group 254: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_983_sample_start_
      -- CP-element group 254: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_980_Update/ack
      -- CP-element group 254: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_980_Update/$exit
      -- CP-element group 254: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_983_Sample/$entry
      -- CP-element group 254: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_983_Sample/req
      -- 
    ack_2024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_980_inst_ack_1, ack => convTranspose_CP_39_elements(254)); -- 
    req_2032_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2032_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(254), ack => WPIPE_Block0_start_983_inst_req_0); -- 
    -- CP-element group 255:  transition  input  output  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	254 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	256 
    -- CP-element group 255:  members (6) 
      -- CP-element group 255: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_983_sample_completed_
      -- CP-element group 255: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_983_update_start_
      -- CP-element group 255: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_983_Sample/$exit
      -- CP-element group 255: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_983_Update/req
      -- CP-element group 255: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_983_Update/$entry
      -- CP-element group 255: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_983_Sample/ack
      -- 
    ack_2033_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_983_inst_ack_0, ack => convTranspose_CP_39_elements(255)); -- 
    req_2037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(255), ack => WPIPE_Block0_start_983_inst_req_1); -- 
    -- CP-element group 256:  transition  input  output  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	255 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	257 
    -- CP-element group 256:  members (6) 
      -- CP-element group 256: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_983_Update/ack
      -- CP-element group 256: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_986_sample_start_
      -- CP-element group 256: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_986_Sample/req
      -- CP-element group 256: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_986_Sample/$entry
      -- CP-element group 256: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_983_update_completed_
      -- CP-element group 256: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_983_Update/$exit
      -- 
    ack_2038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_983_inst_ack_1, ack => convTranspose_CP_39_elements(256)); -- 
    req_2046_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2046_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(256), ack => WPIPE_Block0_start_986_inst_req_0); -- 
    -- CP-element group 257:  transition  input  output  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	256 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	258 
    -- CP-element group 257:  members (6) 
      -- CP-element group 257: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_986_sample_completed_
      -- CP-element group 257: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_986_update_start_
      -- CP-element group 257: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_986_Sample/$exit
      -- CP-element group 257: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_986_Sample/ack
      -- CP-element group 257: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_986_Update/$entry
      -- CP-element group 257: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_986_Update/req
      -- 
    ack_2047_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_986_inst_ack_0, ack => convTranspose_CP_39_elements(257)); -- 
    req_2051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(257), ack => WPIPE_Block0_start_986_inst_req_1); -- 
    -- CP-element group 258:  transition  input  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	257 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	339 
    -- CP-element group 258:  members (3) 
      -- CP-element group 258: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_986_update_completed_
      -- CP-element group 258: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_986_Update/$exit
      -- CP-element group 258: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_986_Update/ack
      -- 
    ack_2052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_986_inst_ack_1, ack => convTranspose_CP_39_elements(258)); -- 
    -- CP-element group 259:  transition  input  output  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	418 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	260 
    -- CP-element group 259:  members (6) 
      -- CP-element group 259: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_989_Update/req
      -- CP-element group 259: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_989_Update/$entry
      -- CP-element group 259: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_989_Sample/ack
      -- CP-element group 259: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_989_Sample/$exit
      -- CP-element group 259: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_989_update_start_
      -- CP-element group 259: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_989_sample_completed_
      -- 
    ack_2061_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_989_inst_ack_0, ack => convTranspose_CP_39_elements(259)); -- 
    req_2065_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2065_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(259), ack => WPIPE_Block1_start_989_inst_req_1); -- 
    -- CP-element group 260:  transition  input  output  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	259 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	261 
    -- CP-element group 260:  members (6) 
      -- CP-element group 260: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_992_Sample/req
      -- CP-element group 260: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_992_Sample/$entry
      -- CP-element group 260: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_992_sample_start_
      -- CP-element group 260: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_989_Update/ack
      -- CP-element group 260: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_989_Update/$exit
      -- CP-element group 260: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_989_update_completed_
      -- 
    ack_2066_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_989_inst_ack_1, ack => convTranspose_CP_39_elements(260)); -- 
    req_2074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(260), ack => WPIPE_Block1_start_992_inst_req_0); -- 
    -- CP-element group 261:  transition  input  output  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	260 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	262 
    -- CP-element group 261:  members (6) 
      -- CP-element group 261: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_992_Sample/$exit
      -- CP-element group 261: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_992_Sample/ack
      -- CP-element group 261: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_992_Update/req
      -- CP-element group 261: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_992_Update/$entry
      -- CP-element group 261: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_992_update_start_
      -- CP-element group 261: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_992_sample_completed_
      -- 
    ack_2075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_992_inst_ack_0, ack => convTranspose_CP_39_elements(261)); -- 
    req_2079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(261), ack => WPIPE_Block1_start_992_inst_req_1); -- 
    -- CP-element group 262:  transition  input  output  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	261 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	263 
    -- CP-element group 262:  members (6) 
      -- CP-element group 262: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_995_Sample/$entry
      -- CP-element group 262: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_992_Update/$exit
      -- CP-element group 262: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_992_Update/ack
      -- CP-element group 262: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_995_sample_start_
      -- CP-element group 262: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_995_Sample/req
      -- CP-element group 262: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_992_update_completed_
      -- 
    ack_2080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_992_inst_ack_1, ack => convTranspose_CP_39_elements(262)); -- 
    req_2088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(262), ack => WPIPE_Block1_start_995_inst_req_0); -- 
    -- CP-element group 263:  transition  input  output  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	262 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	264 
    -- CP-element group 263:  members (6) 
      -- CP-element group 263: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_995_sample_completed_
      -- CP-element group 263: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_995_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_995_Update/req
      -- CP-element group 263: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_995_update_start_
      -- CP-element group 263: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_995_Sample/$exit
      -- CP-element group 263: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_995_Sample/ack
      -- 
    ack_2089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_995_inst_ack_0, ack => convTranspose_CP_39_elements(263)); -- 
    req_2093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(263), ack => WPIPE_Block1_start_995_inst_req_1); -- 
    -- CP-element group 264:  transition  input  output  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	263 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	265 
    -- CP-element group 264:  members (6) 
      -- CP-element group 264: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_995_update_completed_
      -- CP-element group 264: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_995_Update/$exit
      -- CP-element group 264: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_995_Update/ack
      -- CP-element group 264: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_998_sample_start_
      -- CP-element group 264: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_998_Sample/$entry
      -- CP-element group 264: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_998_Sample/req
      -- 
    ack_2094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_995_inst_ack_1, ack => convTranspose_CP_39_elements(264)); -- 
    req_2102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(264), ack => WPIPE_Block1_start_998_inst_req_0); -- 
    -- CP-element group 265:  transition  input  output  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	264 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	266 
    -- CP-element group 265:  members (6) 
      -- CP-element group 265: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_998_sample_completed_
      -- CP-element group 265: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_998_update_start_
      -- CP-element group 265: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_998_Sample/$exit
      -- CP-element group 265: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_998_Sample/ack
      -- CP-element group 265: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_998_Update/$entry
      -- CP-element group 265: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_998_Update/req
      -- 
    ack_2103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_998_inst_ack_0, ack => convTranspose_CP_39_elements(265)); -- 
    req_2107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(265), ack => WPIPE_Block1_start_998_inst_req_1); -- 
    -- CP-element group 266:  transition  input  output  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	265 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	267 
    -- CP-element group 266:  members (6) 
      -- CP-element group 266: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1001_Sample/req
      -- CP-element group 266: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1001_Sample/$entry
      -- CP-element group 266: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_998_update_completed_
      -- CP-element group 266: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_998_Update/$exit
      -- CP-element group 266: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1001_sample_start_
      -- CP-element group 266: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_998_Update/ack
      -- 
    ack_2108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_998_inst_ack_1, ack => convTranspose_CP_39_elements(266)); -- 
    req_2116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(266), ack => WPIPE_Block1_start_1001_inst_req_0); -- 
    -- CP-element group 267:  transition  input  output  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	266 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	268 
    -- CP-element group 267:  members (6) 
      -- CP-element group 267: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1001_sample_completed_
      -- CP-element group 267: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1001_update_start_
      -- CP-element group 267: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1001_Sample/$exit
      -- CP-element group 267: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1001_Sample/ack
      -- CP-element group 267: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1001_Update/$entry
      -- CP-element group 267: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1001_Update/req
      -- 
    ack_2117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1001_inst_ack_0, ack => convTranspose_CP_39_elements(267)); -- 
    req_2121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(267), ack => WPIPE_Block1_start_1001_inst_req_1); -- 
    -- CP-element group 268:  transition  input  output  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	267 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	269 
    -- CP-element group 268:  members (6) 
      -- CP-element group 268: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1001_update_completed_
      -- CP-element group 268: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1001_Update/$exit
      -- CP-element group 268: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1001_Update/ack
      -- CP-element group 268: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1004_Sample/req
      -- CP-element group 268: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1004_Sample/$entry
      -- CP-element group 268: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1004_sample_start_
      -- 
    ack_2122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1001_inst_ack_1, ack => convTranspose_CP_39_elements(268)); -- 
    req_2130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(268), ack => WPIPE_Block1_start_1004_inst_req_0); -- 
    -- CP-element group 269:  transition  input  output  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	268 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	270 
    -- CP-element group 269:  members (6) 
      -- CP-element group 269: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1004_Update/req
      -- CP-element group 269: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1004_Update/$entry
      -- CP-element group 269: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1004_Sample/ack
      -- CP-element group 269: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1004_Sample/$exit
      -- CP-element group 269: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1004_update_start_
      -- CP-element group 269: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1004_sample_completed_
      -- 
    ack_2131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 269_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1004_inst_ack_0, ack => convTranspose_CP_39_elements(269)); -- 
    req_2135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(269), ack => WPIPE_Block1_start_1004_inst_req_1); -- 
    -- CP-element group 270:  transition  input  output  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	269 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	271 
    -- CP-element group 270:  members (6) 
      -- CP-element group 270: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1007_Sample/req
      -- CP-element group 270: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1007_Sample/$entry
      -- CP-element group 270: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1007_sample_start_
      -- CP-element group 270: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1004_Update/ack
      -- CP-element group 270: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1004_Update/$exit
      -- CP-element group 270: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1004_update_completed_
      -- 
    ack_2136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1004_inst_ack_1, ack => convTranspose_CP_39_elements(270)); -- 
    req_2144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(270), ack => WPIPE_Block1_start_1007_inst_req_0); -- 
    -- CP-element group 271:  transition  input  output  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	270 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	272 
    -- CP-element group 271:  members (6) 
      -- CP-element group 271: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1007_Update/req
      -- CP-element group 271: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1007_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1007_Sample/ack
      -- CP-element group 271: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1007_Sample/$exit
      -- CP-element group 271: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1007_update_start_
      -- CP-element group 271: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1007_sample_completed_
      -- 
    ack_2145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1007_inst_ack_0, ack => convTranspose_CP_39_elements(271)); -- 
    req_2149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(271), ack => WPIPE_Block1_start_1007_inst_req_1); -- 
    -- CP-element group 272:  transition  input  output  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	271 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	273 
    -- CP-element group 272:  members (6) 
      -- CP-element group 272: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1010_Sample/req
      -- CP-element group 272: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1010_Sample/$entry
      -- CP-element group 272: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1010_sample_start_
      -- CP-element group 272: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1007_Update/ack
      -- CP-element group 272: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1007_Update/$exit
      -- CP-element group 272: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1007_update_completed_
      -- 
    ack_2150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1007_inst_ack_1, ack => convTranspose_CP_39_elements(272)); -- 
    req_2158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(272), ack => WPIPE_Block1_start_1010_inst_req_0); -- 
    -- CP-element group 273:  transition  input  output  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	272 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	274 
    -- CP-element group 273:  members (6) 
      -- CP-element group 273: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1010_Update/req
      -- CP-element group 273: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1010_Update/$entry
      -- CP-element group 273: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1010_Sample/ack
      -- CP-element group 273: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1010_Sample/$exit
      -- CP-element group 273: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1010_update_start_
      -- CP-element group 273: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1010_sample_completed_
      -- 
    ack_2159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1010_inst_ack_0, ack => convTranspose_CP_39_elements(273)); -- 
    req_2163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(273), ack => WPIPE_Block1_start_1010_inst_req_1); -- 
    -- CP-element group 274:  transition  input  output  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	273 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	275 
    -- CP-element group 274:  members (6) 
      -- CP-element group 274: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1013_Sample/req
      -- CP-element group 274: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1013_Sample/$entry
      -- CP-element group 274: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1013_sample_start_
      -- CP-element group 274: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1010_Update/ack
      -- CP-element group 274: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1010_Update/$exit
      -- CP-element group 274: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1010_update_completed_
      -- 
    ack_2164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1010_inst_ack_1, ack => convTranspose_CP_39_elements(274)); -- 
    req_2172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(274), ack => WPIPE_Block1_start_1013_inst_req_0); -- 
    -- CP-element group 275:  transition  input  output  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	274 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	276 
    -- CP-element group 275:  members (6) 
      -- CP-element group 275: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1013_Update/$entry
      -- CP-element group 275: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1013_Update/req
      -- CP-element group 275: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1013_Sample/ack
      -- CP-element group 275: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1013_Sample/$exit
      -- CP-element group 275: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1013_update_start_
      -- CP-element group 275: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1013_sample_completed_
      -- 
    ack_2173_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1013_inst_ack_0, ack => convTranspose_CP_39_elements(275)); -- 
    req_2177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(275), ack => WPIPE_Block1_start_1013_inst_req_1); -- 
    -- CP-element group 276:  transition  input  output  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	275 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	277 
    -- CP-element group 276:  members (6) 
      -- CP-element group 276: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1013_Update/$exit
      -- CP-element group 276: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1016_Sample/$entry
      -- CP-element group 276: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1013_Update/ack
      -- CP-element group 276: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1016_Sample/req
      -- CP-element group 276: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1016_sample_start_
      -- CP-element group 276: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1013_update_completed_
      -- 
    ack_2178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1013_inst_ack_1, ack => convTranspose_CP_39_elements(276)); -- 
    req_2186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(276), ack => WPIPE_Block1_start_1016_inst_req_0); -- 
    -- CP-element group 277:  transition  input  output  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	276 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	278 
    -- CP-element group 277:  members (6) 
      -- CP-element group 277: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1016_sample_completed_
      -- CP-element group 277: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1016_Update/$entry
      -- CP-element group 277: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1016_Sample/$exit
      -- CP-element group 277: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1016_Update/req
      -- CP-element group 277: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1016_update_start_
      -- CP-element group 277: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1016_Sample/ack
      -- 
    ack_2187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1016_inst_ack_0, ack => convTranspose_CP_39_elements(277)); -- 
    req_2191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(277), ack => WPIPE_Block1_start_1016_inst_req_1); -- 
    -- CP-element group 278:  transition  input  output  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	277 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	279 
    -- CP-element group 278:  members (6) 
      -- CP-element group 278: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1019_sample_start_
      -- CP-element group 278: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1016_update_completed_
      -- CP-element group 278: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1016_Update/$exit
      -- CP-element group 278: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1016_Update/ack
      -- CP-element group 278: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1019_Sample/$entry
      -- CP-element group 278: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1019_Sample/req
      -- 
    ack_2192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1016_inst_ack_1, ack => convTranspose_CP_39_elements(278)); -- 
    req_2200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(278), ack => WPIPE_Block1_start_1019_inst_req_0); -- 
    -- CP-element group 279:  transition  input  output  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	278 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	280 
    -- CP-element group 279:  members (6) 
      -- CP-element group 279: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1019_sample_completed_
      -- CP-element group 279: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1019_update_start_
      -- CP-element group 279: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1019_Update/$entry
      -- CP-element group 279: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1019_Sample/$exit
      -- CP-element group 279: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1019_Sample/ack
      -- CP-element group 279: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1019_Update/req
      -- 
    ack_2201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1019_inst_ack_0, ack => convTranspose_CP_39_elements(279)); -- 
    req_2205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(279), ack => WPIPE_Block1_start_1019_inst_req_1); -- 
    -- CP-element group 280:  transition  input  output  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	279 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	281 
    -- CP-element group 280:  members (6) 
      -- CP-element group 280: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1019_Update/$exit
      -- CP-element group 280: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1019_update_completed_
      -- CP-element group 280: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1019_Update/ack
      -- CP-element group 280: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1022_sample_start_
      -- CP-element group 280: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1022_Sample/$entry
      -- CP-element group 280: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1022_Sample/req
      -- 
    ack_2206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1019_inst_ack_1, ack => convTranspose_CP_39_elements(280)); -- 
    req_2214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(280), ack => WPIPE_Block1_start_1022_inst_req_0); -- 
    -- CP-element group 281:  transition  input  output  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	280 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	282 
    -- CP-element group 281:  members (6) 
      -- CP-element group 281: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1022_sample_completed_
      -- CP-element group 281: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1022_update_start_
      -- CP-element group 281: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1022_Sample/$exit
      -- CP-element group 281: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1022_Sample/ack
      -- CP-element group 281: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1022_Update/$entry
      -- CP-element group 281: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1022_Update/req
      -- 
    ack_2215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1022_inst_ack_0, ack => convTranspose_CP_39_elements(281)); -- 
    req_2219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(281), ack => WPIPE_Block1_start_1022_inst_req_1); -- 
    -- CP-element group 282:  transition  input  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	281 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	339 
    -- CP-element group 282:  members (3) 
      -- CP-element group 282: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1022_update_completed_
      -- CP-element group 282: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1022_Update/ack
      -- CP-element group 282: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1022_Update/$exit
      -- 
    ack_2220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1022_inst_ack_1, ack => convTranspose_CP_39_elements(282)); -- 
    -- CP-element group 283:  transition  input  output  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	418 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	284 
    -- CP-element group 283:  members (6) 
      -- CP-element group 283: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1025_Update/req
      -- CP-element group 283: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1025_Update/$entry
      -- CP-element group 283: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1025_Sample/ack
      -- CP-element group 283: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1025_Sample/$exit
      -- CP-element group 283: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1025_update_start_
      -- CP-element group 283: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1025_sample_completed_
      -- 
    ack_2229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 283_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1025_inst_ack_0, ack => convTranspose_CP_39_elements(283)); -- 
    req_2233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(283), ack => WPIPE_Block2_start_1025_inst_req_1); -- 
    -- CP-element group 284:  transition  input  output  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	283 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	285 
    -- CP-element group 284:  members (6) 
      -- CP-element group 284: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1028_Sample/req
      -- CP-element group 284: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1025_Update/ack
      -- CP-element group 284: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1025_Update/$exit
      -- CP-element group 284: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1028_sample_start_
      -- CP-element group 284: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1028_Sample/$entry
      -- CP-element group 284: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1025_update_completed_
      -- 
    ack_2234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1025_inst_ack_1, ack => convTranspose_CP_39_elements(284)); -- 
    req_2242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(284), ack => WPIPE_Block2_start_1028_inst_req_0); -- 
    -- CP-element group 285:  transition  input  output  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	284 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	286 
    -- CP-element group 285:  members (6) 
      -- CP-element group 285: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1028_Sample/$exit
      -- CP-element group 285: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1028_sample_completed_
      -- CP-element group 285: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1028_update_start_
      -- CP-element group 285: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1028_Sample/ack
      -- CP-element group 285: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1028_Update/$entry
      -- CP-element group 285: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1028_Update/req
      -- 
    ack_2243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1028_inst_ack_0, ack => convTranspose_CP_39_elements(285)); -- 
    req_2247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(285), ack => WPIPE_Block2_start_1028_inst_req_1); -- 
    -- CP-element group 286:  transition  input  output  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	285 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	287 
    -- CP-element group 286:  members (6) 
      -- CP-element group 286: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1028_update_completed_
      -- CP-element group 286: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1028_Update/$exit
      -- CP-element group 286: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1031_Sample/req
      -- CP-element group 286: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1031_Sample/$entry
      -- CP-element group 286: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1031_sample_start_
      -- CP-element group 286: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1028_Update/ack
      -- 
    ack_2248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1028_inst_ack_1, ack => convTranspose_CP_39_elements(286)); -- 
    req_2256_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2256_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(286), ack => WPIPE_Block2_start_1031_inst_req_0); -- 
    -- CP-element group 287:  transition  input  output  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	286 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	288 
    -- CP-element group 287:  members (6) 
      -- CP-element group 287: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1031_Update/req
      -- CP-element group 287: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1031_Update/$entry
      -- CP-element group 287: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1031_Sample/ack
      -- CP-element group 287: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1031_Sample/$exit
      -- CP-element group 287: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1031_update_start_
      -- CP-element group 287: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1031_sample_completed_
      -- 
    ack_2257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1031_inst_ack_0, ack => convTranspose_CP_39_elements(287)); -- 
    req_2261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(287), ack => WPIPE_Block2_start_1031_inst_req_1); -- 
    -- CP-element group 288:  transition  input  output  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	287 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	289 
    -- CP-element group 288:  members (6) 
      -- CP-element group 288: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1034_Sample/req
      -- CP-element group 288: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1034_Sample/$entry
      -- CP-element group 288: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1034_sample_start_
      -- CP-element group 288: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1031_Update/ack
      -- CP-element group 288: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1031_Update/$exit
      -- CP-element group 288: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1031_update_completed_
      -- 
    ack_2262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1031_inst_ack_1, ack => convTranspose_CP_39_elements(288)); -- 
    req_2270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(288), ack => WPIPE_Block2_start_1034_inst_req_0); -- 
    -- CP-element group 289:  transition  input  output  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	288 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	290 
    -- CP-element group 289:  members (6) 
      -- CP-element group 289: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1034_Update/req
      -- CP-element group 289: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1034_Update/$entry
      -- CP-element group 289: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1034_Sample/ack
      -- CP-element group 289: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1034_Sample/$exit
      -- CP-element group 289: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1034_update_start_
      -- CP-element group 289: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1034_sample_completed_
      -- 
    ack_2271_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1034_inst_ack_0, ack => convTranspose_CP_39_elements(289)); -- 
    req_2275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(289), ack => WPIPE_Block2_start_1034_inst_req_1); -- 
    -- CP-element group 290:  transition  input  output  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	289 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	291 
    -- CP-element group 290:  members (6) 
      -- CP-element group 290: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1037_Sample/req
      -- CP-element group 290: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1037_Sample/$entry
      -- CP-element group 290: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1037_sample_start_
      -- CP-element group 290: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1034_Update/ack
      -- CP-element group 290: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1034_Update/$exit
      -- CP-element group 290: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1034_update_completed_
      -- 
    ack_2276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1034_inst_ack_1, ack => convTranspose_CP_39_elements(290)); -- 
    req_2284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(290), ack => WPIPE_Block2_start_1037_inst_req_0); -- 
    -- CP-element group 291:  transition  input  output  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	290 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	292 
    -- CP-element group 291:  members (6) 
      -- CP-element group 291: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1037_Update/$entry
      -- CP-element group 291: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1037_Sample/ack
      -- CP-element group 291: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1037_Update/req
      -- CP-element group 291: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1037_Sample/$exit
      -- CP-element group 291: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1037_update_start_
      -- CP-element group 291: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1037_sample_completed_
      -- 
    ack_2285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1037_inst_ack_0, ack => convTranspose_CP_39_elements(291)); -- 
    req_2289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(291), ack => WPIPE_Block2_start_1037_inst_req_1); -- 
    -- CP-element group 292:  transition  input  output  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	291 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	293 
    -- CP-element group 292:  members (6) 
      -- CP-element group 292: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1037_Update/ack
      -- CP-element group 292: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1037_Update/$exit
      -- CP-element group 292: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1040_Sample/$entry
      -- CP-element group 292: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1040_Sample/req
      -- CP-element group 292: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1040_sample_start_
      -- CP-element group 292: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1037_update_completed_
      -- 
    ack_2290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1037_inst_ack_1, ack => convTranspose_CP_39_elements(292)); -- 
    req_2298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(292), ack => WPIPE_Block2_start_1040_inst_req_0); -- 
    -- CP-element group 293:  transition  input  output  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	292 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	294 
    -- CP-element group 293:  members (6) 
      -- CP-element group 293: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1040_sample_completed_
      -- CP-element group 293: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1040_Sample/$exit
      -- CP-element group 293: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1040_Sample/ack
      -- CP-element group 293: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1040_update_start_
      -- CP-element group 293: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1040_Update/$entry
      -- CP-element group 293: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1040_Update/req
      -- 
    ack_2299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 293_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1040_inst_ack_0, ack => convTranspose_CP_39_elements(293)); -- 
    req_2303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(293), ack => WPIPE_Block2_start_1040_inst_req_1); -- 
    -- CP-element group 294:  transition  input  output  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	293 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	295 
    -- CP-element group 294:  members (6) 
      -- CP-element group 294: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1040_Update/$exit
      -- CP-element group 294: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1043_Sample/req
      -- CP-element group 294: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1040_Update/ack
      -- CP-element group 294: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1043_sample_start_
      -- CP-element group 294: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1040_update_completed_
      -- CP-element group 294: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1043_Sample/$entry
      -- 
    ack_2304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 294_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1040_inst_ack_1, ack => convTranspose_CP_39_elements(294)); -- 
    req_2312_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2312_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(294), ack => WPIPE_Block2_start_1043_inst_req_0); -- 
    -- CP-element group 295:  transition  input  output  bypass 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	294 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	296 
    -- CP-element group 295:  members (6) 
      -- CP-element group 295: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1043_Update/req
      -- CP-element group 295: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1043_sample_completed_
      -- CP-element group 295: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1043_update_start_
      -- CP-element group 295: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1043_Sample/$exit
      -- CP-element group 295: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1043_Sample/ack
      -- CP-element group 295: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1043_Update/$entry
      -- 
    ack_2313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1043_inst_ack_0, ack => convTranspose_CP_39_elements(295)); -- 
    req_2317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(295), ack => WPIPE_Block2_start_1043_inst_req_1); -- 
    -- CP-element group 296:  transition  input  output  bypass 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	295 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	297 
    -- CP-element group 296:  members (6) 
      -- CP-element group 296: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1043_update_completed_
      -- CP-element group 296: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1043_Update/$exit
      -- CP-element group 296: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1046_Sample/req
      -- CP-element group 296: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1046_Sample/$entry
      -- CP-element group 296: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1046_sample_start_
      -- CP-element group 296: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1043_Update/ack
      -- 
    ack_2318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1043_inst_ack_1, ack => convTranspose_CP_39_elements(296)); -- 
    req_2326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(296), ack => WPIPE_Block2_start_1046_inst_req_0); -- 
    -- CP-element group 297:  transition  input  output  bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	296 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	298 
    -- CP-element group 297:  members (6) 
      -- CP-element group 297: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1046_Update/$entry
      -- CP-element group 297: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1046_Update/req
      -- CP-element group 297: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1046_Sample/ack
      -- CP-element group 297: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1046_Sample/$exit
      -- CP-element group 297: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1046_update_start_
      -- CP-element group 297: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1046_sample_completed_
      -- 
    ack_2327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1046_inst_ack_0, ack => convTranspose_CP_39_elements(297)); -- 
    req_2331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(297), ack => WPIPE_Block2_start_1046_inst_req_1); -- 
    -- CP-element group 298:  transition  input  output  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	297 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	299 
    -- CP-element group 298:  members (6) 
      -- CP-element group 298: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1046_Update/$exit
      -- CP-element group 298: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1046_Update/ack
      -- CP-element group 298: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1049_sample_start_
      -- CP-element group 298: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1049_Sample/$entry
      -- CP-element group 298: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1049_Sample/req
      -- CP-element group 298: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1046_update_completed_
      -- 
    ack_2332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 298_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1046_inst_ack_1, ack => convTranspose_CP_39_elements(298)); -- 
    req_2340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(298), ack => WPIPE_Block2_start_1049_inst_req_0); -- 
    -- CP-element group 299:  transition  input  output  bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	298 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	300 
    -- CP-element group 299:  members (6) 
      -- CP-element group 299: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1049_sample_completed_
      -- CP-element group 299: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1049_update_start_
      -- CP-element group 299: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1049_Sample/$exit
      -- CP-element group 299: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1049_Update/req
      -- CP-element group 299: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1049_Update/$entry
      -- CP-element group 299: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1049_Sample/ack
      -- 
    ack_2341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1049_inst_ack_0, ack => convTranspose_CP_39_elements(299)); -- 
    req_2345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(299), ack => WPIPE_Block2_start_1049_inst_req_1); -- 
    -- CP-element group 300:  transition  input  output  bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	299 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	301 
    -- CP-element group 300:  members (6) 
      -- CP-element group 300: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1052_sample_start_
      -- CP-element group 300: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1049_update_completed_
      -- CP-element group 300: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1049_Update/ack
      -- CP-element group 300: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1049_Update/$exit
      -- CP-element group 300: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1052_Sample/req
      -- CP-element group 300: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1052_Sample/$entry
      -- 
    ack_2346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1049_inst_ack_1, ack => convTranspose_CP_39_elements(300)); -- 
    req_2354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(300), ack => WPIPE_Block2_start_1052_inst_req_0); -- 
    -- CP-element group 301:  transition  input  output  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	300 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	302 
    -- CP-element group 301:  members (6) 
      -- CP-element group 301: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1052_Update/req
      -- CP-element group 301: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1052_sample_completed_
      -- CP-element group 301: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1052_update_start_
      -- CP-element group 301: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1052_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1052_Sample/ack
      -- CP-element group 301: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1052_Sample/$exit
      -- 
    ack_2355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 301_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1052_inst_ack_0, ack => convTranspose_CP_39_elements(301)); -- 
    req_2359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(301), ack => WPIPE_Block2_start_1052_inst_req_1); -- 
    -- CP-element group 302:  transition  input  output  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	301 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	303 
    -- CP-element group 302:  members (6) 
      -- CP-element group 302: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1052_Update/ack
      -- CP-element group 302: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1052_update_completed_
      -- CP-element group 302: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1052_Update/$exit
      -- CP-element group 302: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1055_Sample/req
      -- CP-element group 302: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1055_Sample/$entry
      -- CP-element group 302: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1055_sample_start_
      -- 
    ack_2360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 302_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1052_inst_ack_1, ack => convTranspose_CP_39_elements(302)); -- 
    req_2368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(302), ack => WPIPE_Block2_start_1055_inst_req_0); -- 
    -- CP-element group 303:  transition  input  output  bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	302 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	304 
    -- CP-element group 303:  members (6) 
      -- CP-element group 303: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1055_Update/req
      -- CP-element group 303: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1055_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1055_Sample/ack
      -- CP-element group 303: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1055_Sample/$exit
      -- CP-element group 303: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1055_update_start_
      -- CP-element group 303: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1055_sample_completed_
      -- 
    ack_2369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1055_inst_ack_0, ack => convTranspose_CP_39_elements(303)); -- 
    req_2373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(303), ack => WPIPE_Block2_start_1055_inst_req_1); -- 
    -- CP-element group 304:  transition  input  output  bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	303 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	305 
    -- CP-element group 304:  members (6) 
      -- CP-element group 304: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1055_Update/ack
      -- CP-element group 304: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1055_Update/$exit
      -- CP-element group 304: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1058_Sample/req
      -- CP-element group 304: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1058_Sample/$entry
      -- CP-element group 304: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1055_update_completed_
      -- CP-element group 304: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1058_sample_start_
      -- 
    ack_2374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1055_inst_ack_1, ack => convTranspose_CP_39_elements(304)); -- 
    req_2382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(304), ack => WPIPE_Block2_start_1058_inst_req_0); -- 
    -- CP-element group 305:  transition  input  output  bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	304 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	306 
    -- CP-element group 305:  members (6) 
      -- CP-element group 305: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1058_Update/req
      -- CP-element group 305: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1058_Update/$entry
      -- CP-element group 305: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1058_Sample/ack
      -- CP-element group 305: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1058_Sample/$exit
      -- CP-element group 305: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1058_update_start_
      -- CP-element group 305: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1058_sample_completed_
      -- 
    ack_2383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 305_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1058_inst_ack_0, ack => convTranspose_CP_39_elements(305)); -- 
    req_2387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(305), ack => WPIPE_Block2_start_1058_inst_req_1); -- 
    -- CP-element group 306:  transition  input  bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	305 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	339 
    -- CP-element group 306:  members (3) 
      -- CP-element group 306: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1058_Update/ack
      -- CP-element group 306: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1058_Update/$exit
      -- CP-element group 306: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1058_update_completed_
      -- 
    ack_2388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1058_inst_ack_1, ack => convTranspose_CP_39_elements(306)); -- 
    -- CP-element group 307:  transition  input  output  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	418 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	308 
    -- CP-element group 307:  members (6) 
      -- CP-element group 307: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1061_Sample/ack
      -- CP-element group 307: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1061_Update/$entry
      -- CP-element group 307: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1061_Update/req
      -- CP-element group 307: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1061_Sample/$exit
      -- CP-element group 307: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1061_update_start_
      -- CP-element group 307: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1061_sample_completed_
      -- 
    ack_2397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1061_inst_ack_0, ack => convTranspose_CP_39_elements(307)); -- 
    req_2401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(307), ack => WPIPE_Block3_start_1061_inst_req_1); -- 
    -- CP-element group 308:  transition  input  output  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	307 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	309 
    -- CP-element group 308:  members (6) 
      -- CP-element group 308: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1061_Update/$exit
      -- CP-element group 308: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1064_Sample/$entry
      -- CP-element group 308: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1061_Update/ack
      -- CP-element group 308: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1064_Sample/req
      -- CP-element group 308: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1064_sample_start_
      -- CP-element group 308: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1061_update_completed_
      -- 
    ack_2402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1061_inst_ack_1, ack => convTranspose_CP_39_elements(308)); -- 
    req_2410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(308), ack => WPIPE_Block3_start_1064_inst_req_0); -- 
    -- CP-element group 309:  transition  input  output  bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	308 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	310 
    -- CP-element group 309:  members (6) 
      -- CP-element group 309: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1064_update_start_
      -- CP-element group 309: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1064_sample_completed_
      -- CP-element group 309: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1064_Sample/$exit
      -- CP-element group 309: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1064_Update/req
      -- CP-element group 309: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1064_Update/$entry
      -- CP-element group 309: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1064_Sample/ack
      -- 
    ack_2411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 309_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1064_inst_ack_0, ack => convTranspose_CP_39_elements(309)); -- 
    req_2415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(309), ack => WPIPE_Block3_start_1064_inst_req_1); -- 
    -- CP-element group 310:  transition  input  output  bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	309 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	311 
    -- CP-element group 310:  members (6) 
      -- CP-element group 310: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1067_Sample/$entry
      -- CP-element group 310: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1064_update_completed_
      -- CP-element group 310: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1067_Sample/req
      -- CP-element group 310: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1067_sample_start_
      -- CP-element group 310: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1064_Update/ack
      -- CP-element group 310: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1064_Update/$exit
      -- 
    ack_2416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 310_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1064_inst_ack_1, ack => convTranspose_CP_39_elements(310)); -- 
    req_2424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(310), ack => WPIPE_Block3_start_1067_inst_req_0); -- 
    -- CP-element group 311:  transition  input  output  bypass 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	310 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	312 
    -- CP-element group 311:  members (6) 
      -- CP-element group 311: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1067_Sample/ack
      -- CP-element group 311: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1067_Sample/$exit
      -- CP-element group 311: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1067_sample_completed_
      -- CP-element group 311: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1067_Update/req
      -- CP-element group 311: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1067_Update/$entry
      -- CP-element group 311: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1067_update_start_
      -- 
    ack_2425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1067_inst_ack_0, ack => convTranspose_CP_39_elements(311)); -- 
    req_2429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(311), ack => WPIPE_Block3_start_1067_inst_req_1); -- 
    -- CP-element group 312:  transition  input  output  bypass 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	311 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	313 
    -- CP-element group 312:  members (6) 
      -- CP-element group 312: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1067_update_completed_
      -- CP-element group 312: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1067_Update/ack
      -- CP-element group 312: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1067_Update/$exit
      -- CP-element group 312: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1070_sample_start_
      -- CP-element group 312: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1070_Sample/$entry
      -- CP-element group 312: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1070_Sample/req
      -- 
    ack_2430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1067_inst_ack_1, ack => convTranspose_CP_39_elements(312)); -- 
    req_2438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(312), ack => WPIPE_Block3_start_1070_inst_req_0); -- 
    -- CP-element group 313:  transition  input  output  bypass 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	312 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	314 
    -- CP-element group 313:  members (6) 
      -- CP-element group 313: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1070_sample_completed_
      -- CP-element group 313: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1070_update_start_
      -- CP-element group 313: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1070_Sample/$exit
      -- CP-element group 313: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1070_Sample/ack
      -- CP-element group 313: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1070_Update/$entry
      -- CP-element group 313: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1070_Update/req
      -- 
    ack_2439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1070_inst_ack_0, ack => convTranspose_CP_39_elements(313)); -- 
    req_2443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(313), ack => WPIPE_Block3_start_1070_inst_req_1); -- 
    -- CP-element group 314:  transition  input  output  bypass 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	313 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	315 
    -- CP-element group 314:  members (6) 
      -- CP-element group 314: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1070_update_completed_
      -- CP-element group 314: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1070_Update/$exit
      -- CP-element group 314: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1070_Update/ack
      -- CP-element group 314: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1073_sample_start_
      -- CP-element group 314: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1073_Sample/$entry
      -- CP-element group 314: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1073_Sample/req
      -- 
    ack_2444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1070_inst_ack_1, ack => convTranspose_CP_39_elements(314)); -- 
    req_2452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(314), ack => WPIPE_Block3_start_1073_inst_req_0); -- 
    -- CP-element group 315:  transition  input  output  bypass 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	314 
    -- CP-element group 315: successors 
    -- CP-element group 315: 	316 
    -- CP-element group 315:  members (6) 
      -- CP-element group 315: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1073_Update/$entry
      -- CP-element group 315: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1073_sample_completed_
      -- CP-element group 315: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1073_update_start_
      -- CP-element group 315: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1073_Sample/$exit
      -- CP-element group 315: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1073_Sample/ack
      -- CP-element group 315: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1073_Update/req
      -- 
    ack_2453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1073_inst_ack_0, ack => convTranspose_CP_39_elements(315)); -- 
    req_2457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(315), ack => WPIPE_Block3_start_1073_inst_req_1); -- 
    -- CP-element group 316:  transition  input  output  bypass 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	315 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	317 
    -- CP-element group 316:  members (6) 
      -- CP-element group 316: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1073_Update/$exit
      -- CP-element group 316: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1073_update_completed_
      -- CP-element group 316: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1073_Update/ack
      -- CP-element group 316: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1076_sample_start_
      -- CP-element group 316: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1076_Sample/$entry
      -- CP-element group 316: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1076_Sample/req
      -- 
    ack_2458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1073_inst_ack_1, ack => convTranspose_CP_39_elements(316)); -- 
    req_2466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(316), ack => WPIPE_Block3_start_1076_inst_req_0); -- 
    -- CP-element group 317:  transition  input  output  bypass 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	316 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	318 
    -- CP-element group 317:  members (6) 
      -- CP-element group 317: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1076_sample_completed_
      -- CP-element group 317: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1076_update_start_
      -- CP-element group 317: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1076_Sample/$exit
      -- CP-element group 317: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1076_Sample/ack
      -- CP-element group 317: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1076_Update/$entry
      -- CP-element group 317: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1076_Update/req
      -- 
    ack_2467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 317_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1076_inst_ack_0, ack => convTranspose_CP_39_elements(317)); -- 
    req_2471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(317), ack => WPIPE_Block3_start_1076_inst_req_1); -- 
    -- CP-element group 318:  transition  input  output  bypass 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	317 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	319 
    -- CP-element group 318:  members (6) 
      -- CP-element group 318: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1076_update_completed_
      -- CP-element group 318: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1076_Update/$exit
      -- CP-element group 318: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1076_Update/ack
      -- CP-element group 318: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1079_sample_start_
      -- CP-element group 318: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1079_Sample/$entry
      -- CP-element group 318: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1079_Sample/req
      -- 
    ack_2472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 318_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1076_inst_ack_1, ack => convTranspose_CP_39_elements(318)); -- 
    req_2480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(318), ack => WPIPE_Block3_start_1079_inst_req_0); -- 
    -- CP-element group 319:  transition  input  output  bypass 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	318 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	320 
    -- CP-element group 319:  members (6) 
      -- CP-element group 319: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1079_sample_completed_
      -- CP-element group 319: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1079_update_start_
      -- CP-element group 319: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1079_Sample/$exit
      -- CP-element group 319: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1079_Sample/ack
      -- CP-element group 319: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1079_Update/$entry
      -- CP-element group 319: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1079_Update/req
      -- 
    ack_2481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 319_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1079_inst_ack_0, ack => convTranspose_CP_39_elements(319)); -- 
    req_2485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(319), ack => WPIPE_Block3_start_1079_inst_req_1); -- 
    -- CP-element group 320:  transition  input  output  bypass 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	319 
    -- CP-element group 320: successors 
    -- CP-element group 320: 	321 
    -- CP-element group 320:  members (6) 
      -- CP-element group 320: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1079_update_completed_
      -- CP-element group 320: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1079_Update/$exit
      -- CP-element group 320: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1079_Update/ack
      -- CP-element group 320: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1082_sample_start_
      -- CP-element group 320: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1082_Sample/$entry
      -- CP-element group 320: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1082_Sample/req
      -- 
    ack_2486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 320_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1079_inst_ack_1, ack => convTranspose_CP_39_elements(320)); -- 
    req_2494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(320), ack => WPIPE_Block3_start_1082_inst_req_0); -- 
    -- CP-element group 321:  transition  input  output  bypass 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	320 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	322 
    -- CP-element group 321:  members (6) 
      -- CP-element group 321: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1082_sample_completed_
      -- CP-element group 321: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1082_update_start_
      -- CP-element group 321: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1082_Sample/$exit
      -- CP-element group 321: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1082_Sample/ack
      -- CP-element group 321: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1082_Update/$entry
      -- CP-element group 321: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1082_Update/req
      -- 
    ack_2495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1082_inst_ack_0, ack => convTranspose_CP_39_elements(321)); -- 
    req_2499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(321), ack => WPIPE_Block3_start_1082_inst_req_1); -- 
    -- CP-element group 322:  transition  input  output  bypass 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	321 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	323 
    -- CP-element group 322:  members (6) 
      -- CP-element group 322: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1082_update_completed_
      -- CP-element group 322: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1082_Update/$exit
      -- CP-element group 322: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1082_Update/ack
      -- CP-element group 322: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1085_sample_start_
      -- CP-element group 322: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1085_Sample/$entry
      -- CP-element group 322: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1085_Sample/req
      -- 
    ack_2500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 322_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1082_inst_ack_1, ack => convTranspose_CP_39_elements(322)); -- 
    req_2508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(322), ack => WPIPE_Block3_start_1085_inst_req_0); -- 
    -- CP-element group 323:  transition  input  output  bypass 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	322 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	324 
    -- CP-element group 323:  members (6) 
      -- CP-element group 323: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1085_sample_completed_
      -- CP-element group 323: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1085_update_start_
      -- CP-element group 323: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1085_Sample/$exit
      -- CP-element group 323: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1085_Sample/ack
      -- CP-element group 323: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1085_Update/$entry
      -- CP-element group 323: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1085_Update/req
      -- 
    ack_2509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 323_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1085_inst_ack_0, ack => convTranspose_CP_39_elements(323)); -- 
    req_2513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(323), ack => WPIPE_Block3_start_1085_inst_req_1); -- 
    -- CP-element group 324:  transition  input  output  bypass 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	323 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	325 
    -- CP-element group 324:  members (6) 
      -- CP-element group 324: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1085_update_completed_
      -- CP-element group 324: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1085_Update/$exit
      -- CP-element group 324: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1085_Update/ack
      -- CP-element group 324: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1088_sample_start_
      -- CP-element group 324: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1088_Sample/$entry
      -- CP-element group 324: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1088_Sample/req
      -- 
    ack_2514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 324_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1085_inst_ack_1, ack => convTranspose_CP_39_elements(324)); -- 
    req_2522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(324), ack => WPIPE_Block3_start_1088_inst_req_0); -- 
    -- CP-element group 325:  transition  input  output  bypass 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	324 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	326 
    -- CP-element group 325:  members (6) 
      -- CP-element group 325: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1088_sample_completed_
      -- CP-element group 325: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1088_update_start_
      -- CP-element group 325: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1088_Sample/$exit
      -- CP-element group 325: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1088_Sample/ack
      -- CP-element group 325: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1088_Update/$entry
      -- CP-element group 325: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1088_Update/req
      -- 
    ack_2523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 325_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1088_inst_ack_0, ack => convTranspose_CP_39_elements(325)); -- 
    req_2527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(325), ack => WPIPE_Block3_start_1088_inst_req_1); -- 
    -- CP-element group 326:  transition  input  output  bypass 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	325 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	327 
    -- CP-element group 326:  members (6) 
      -- CP-element group 326: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1088_update_completed_
      -- CP-element group 326: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1088_Update/$exit
      -- CP-element group 326: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1088_Update/ack
      -- CP-element group 326: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1091_sample_start_
      -- CP-element group 326: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1091_Sample/$entry
      -- CP-element group 326: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1091_Sample/req
      -- 
    ack_2528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 326_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1088_inst_ack_1, ack => convTranspose_CP_39_elements(326)); -- 
    req_2536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(326), ack => WPIPE_Block3_start_1091_inst_req_0); -- 
    -- CP-element group 327:  transition  input  output  bypass 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	326 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	328 
    -- CP-element group 327:  members (6) 
      -- CP-element group 327: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1091_sample_completed_
      -- CP-element group 327: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1091_update_start_
      -- CP-element group 327: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1091_Sample/$exit
      -- CP-element group 327: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1091_Sample/ack
      -- CP-element group 327: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1091_Update/$entry
      -- CP-element group 327: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1091_Update/req
      -- 
    ack_2537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 327_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1091_inst_ack_0, ack => convTranspose_CP_39_elements(327)); -- 
    req_2541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(327), ack => WPIPE_Block3_start_1091_inst_req_1); -- 
    -- CP-element group 328:  transition  input  output  bypass 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	327 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	329 
    -- CP-element group 328:  members (6) 
      -- CP-element group 328: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1091_update_completed_
      -- CP-element group 328: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1091_Update/$exit
      -- CP-element group 328: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1091_Update/ack
      -- CP-element group 328: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1094_sample_start_
      -- CP-element group 328: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1094_Sample/$entry
      -- CP-element group 328: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1094_Sample/req
      -- 
    ack_2542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 328_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1091_inst_ack_1, ack => convTranspose_CP_39_elements(328)); -- 
    req_2550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(328), ack => WPIPE_Block3_start_1094_inst_req_0); -- 
    -- CP-element group 329:  transition  input  output  bypass 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	328 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	330 
    -- CP-element group 329:  members (6) 
      -- CP-element group 329: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1094_sample_completed_
      -- CP-element group 329: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1094_update_start_
      -- CP-element group 329: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1094_Sample/$exit
      -- CP-element group 329: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1094_Sample/ack
      -- CP-element group 329: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1094_Update/$entry
      -- CP-element group 329: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1094_Update/req
      -- 
    ack_2551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 329_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1094_inst_ack_0, ack => convTranspose_CP_39_elements(329)); -- 
    req_2555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(329), ack => WPIPE_Block3_start_1094_inst_req_1); -- 
    -- CP-element group 330:  transition  input  bypass 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	329 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	339 
    -- CP-element group 330:  members (3) 
      -- CP-element group 330: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1094_update_completed_
      -- CP-element group 330: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1094_Update/$exit
      -- CP-element group 330: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1094_Update/ack
      -- 
    ack_2556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 330_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1094_inst_ack_1, ack => convTranspose_CP_39_elements(330)); -- 
    -- CP-element group 331:  transition  input  output  bypass 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	418 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	332 
    -- CP-element group 331:  members (6) 
      -- CP-element group 331: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block0_done_1098_sample_completed_
      -- CP-element group 331: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block0_done_1098_update_start_
      -- CP-element group 331: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block0_done_1098_Sample/$exit
      -- CP-element group 331: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block0_done_1098_Sample/ra
      -- CP-element group 331: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block0_done_1098_Update/$entry
      -- CP-element group 331: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block0_done_1098_Update/cr
      -- 
    ra_2565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 331_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1098_inst_ack_0, ack => convTranspose_CP_39_elements(331)); -- 
    cr_2569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(331), ack => RPIPE_Block0_done_1098_inst_req_1); -- 
    -- CP-element group 332:  transition  input  bypass 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	331 
    -- CP-element group 332: successors 
    -- CP-element group 332: 	339 
    -- CP-element group 332:  members (3) 
      -- CP-element group 332: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block0_done_1098_update_completed_
      -- CP-element group 332: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block0_done_1098_Update/$exit
      -- CP-element group 332: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block0_done_1098_Update/ca
      -- 
    ca_2570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1098_inst_ack_1, ack => convTranspose_CP_39_elements(332)); -- 
    -- CP-element group 333:  transition  input  output  bypass 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	418 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	334 
    -- CP-element group 333:  members (6) 
      -- CP-element group 333: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block1_done_1101_sample_completed_
      -- CP-element group 333: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block1_done_1101_update_start_
      -- CP-element group 333: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block1_done_1101_Sample/$exit
      -- CP-element group 333: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block1_done_1101_Sample/ra
      -- CP-element group 333: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block1_done_1101_Update/$entry
      -- CP-element group 333: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block1_done_1101_Update/cr
      -- 
    ra_2579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 333_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1101_inst_ack_0, ack => convTranspose_CP_39_elements(333)); -- 
    cr_2583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(333), ack => RPIPE_Block1_done_1101_inst_req_1); -- 
    -- CP-element group 334:  transition  input  bypass 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	333 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	339 
    -- CP-element group 334:  members (3) 
      -- CP-element group 334: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block1_done_1101_update_completed_
      -- CP-element group 334: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block1_done_1101_Update/$exit
      -- CP-element group 334: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block1_done_1101_Update/ca
      -- 
    ca_2584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 334_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1101_inst_ack_1, ack => convTranspose_CP_39_elements(334)); -- 
    -- CP-element group 335:  transition  input  output  bypass 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	418 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	336 
    -- CP-element group 335:  members (6) 
      -- CP-element group 335: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block2_done_1104_sample_completed_
      -- CP-element group 335: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block2_done_1104_update_start_
      -- CP-element group 335: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block2_done_1104_Sample/$exit
      -- CP-element group 335: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block2_done_1104_Sample/ra
      -- CP-element group 335: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block2_done_1104_Update/$entry
      -- CP-element group 335: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block2_done_1104_Update/cr
      -- 
    ra_2593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 335_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1104_inst_ack_0, ack => convTranspose_CP_39_elements(335)); -- 
    cr_2597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(335), ack => RPIPE_Block2_done_1104_inst_req_1); -- 
    -- CP-element group 336:  transition  input  bypass 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	335 
    -- CP-element group 336: successors 
    -- CP-element group 336: 	339 
    -- CP-element group 336:  members (3) 
      -- CP-element group 336: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block2_done_1104_update_completed_
      -- CP-element group 336: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block2_done_1104_Update/$exit
      -- CP-element group 336: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block2_done_1104_Update/ca
      -- 
    ca_2598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1104_inst_ack_1, ack => convTranspose_CP_39_elements(336)); -- 
    -- CP-element group 337:  transition  input  output  bypass 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	418 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	338 
    -- CP-element group 337:  members (6) 
      -- CP-element group 337: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block3_done_1107_sample_completed_
      -- CP-element group 337: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block3_done_1107_update_start_
      -- CP-element group 337: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block3_done_1107_Sample/$exit
      -- CP-element group 337: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block3_done_1107_Sample/ra
      -- CP-element group 337: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block3_done_1107_Update/$entry
      -- CP-element group 337: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block3_done_1107_Update/cr
      -- 
    ra_2607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1107_inst_ack_0, ack => convTranspose_CP_39_elements(337)); -- 
    cr_2611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(337), ack => RPIPE_Block3_done_1107_inst_req_1); -- 
    -- CP-element group 338:  transition  input  bypass 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	337 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	339 
    -- CP-element group 338:  members (3) 
      -- CP-element group 338: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block3_done_1107_update_completed_
      -- CP-element group 338: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block3_done_1107_Update/$exit
      -- CP-element group 338: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block3_done_1107_Update/ca
      -- 
    ca_2612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 338_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1107_inst_ack_1, ack => convTranspose_CP_39_elements(338)); -- 
    -- CP-element group 339:  join  fork  transition  place  output  bypass 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	282 
    -- CP-element group 339: 	306 
    -- CP-element group 339: 	330 
    -- CP-element group 339: 	332 
    -- CP-element group 339: 	334 
    -- CP-element group 339: 	336 
    -- CP-element group 339: 	338 
    -- CP-element group 339: 	234 
    -- CP-element group 339: 	258 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	340 
    -- CP-element group 339: 	341 
    -- CP-element group 339: 	343 
    -- CP-element group 339:  members (13) 
      -- CP-element group 339: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108__exit__
      -- CP-element group 339: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124__entry__
      -- CP-element group 339: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/$exit
      -- CP-element group 339: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/$entry
      -- CP-element group 339: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/call_stmt_1111_sample_start_
      -- CP-element group 339: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/call_stmt_1111_update_start_
      -- CP-element group 339: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/call_stmt_1111_Sample/$entry
      -- CP-element group 339: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/call_stmt_1111_Sample/crr
      -- CP-element group 339: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/call_stmt_1111_Update/$entry
      -- CP-element group 339: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/call_stmt_1111_Update/ccr
      -- CP-element group 339: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/type_cast_1115_update_start_
      -- CP-element group 339: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/type_cast_1115_Update/$entry
      -- CP-element group 339: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/type_cast_1115_Update/cr
      -- 
    crr_2623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(339), ack => call_stmt_1111_call_req_0); -- 
    ccr_2628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(339), ack => call_stmt_1111_call_req_1); -- 
    cr_2642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(339), ack => type_cast_1115_inst_req_1); -- 
    convTranspose_cp_element_group_339: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_339"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(282) & convTranspose_CP_39_elements(306) & convTranspose_CP_39_elements(330) & convTranspose_CP_39_elements(332) & convTranspose_CP_39_elements(334) & convTranspose_CP_39_elements(336) & convTranspose_CP_39_elements(338) & convTranspose_CP_39_elements(234) & convTranspose_CP_39_elements(258);
      gj_convTranspose_cp_element_group_339 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(339), clk => clk, reset => reset); --
    end block;
    -- CP-element group 340:  transition  input  bypass 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	339 
    -- CP-element group 340: successors 
    -- CP-element group 340:  members (3) 
      -- CP-element group 340: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/call_stmt_1111_sample_completed_
      -- CP-element group 340: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/call_stmt_1111_Sample/$exit
      -- CP-element group 340: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/call_stmt_1111_Sample/cra
      -- 
    cra_2624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1111_call_ack_0, ack => convTranspose_CP_39_elements(340)); -- 
    -- CP-element group 341:  transition  input  output  bypass 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	339 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	342 
    -- CP-element group 341:  members (6) 
      -- CP-element group 341: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/call_stmt_1111_update_completed_
      -- CP-element group 341: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/call_stmt_1111_Update/$exit
      -- CP-element group 341: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/call_stmt_1111_Update/cca
      -- CP-element group 341: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/type_cast_1115_sample_start_
      -- CP-element group 341: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/type_cast_1115_Sample/$entry
      -- CP-element group 341: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/type_cast_1115_Sample/rr
      -- 
    cca_2629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1111_call_ack_1, ack => convTranspose_CP_39_elements(341)); -- 
    rr_2637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(341), ack => type_cast_1115_inst_req_0); -- 
    -- CP-element group 342:  transition  input  bypass 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	341 
    -- CP-element group 342: successors 
    -- CP-element group 342:  members (3) 
      -- CP-element group 342: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/type_cast_1115_sample_completed_
      -- CP-element group 342: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/type_cast_1115_Sample/$exit
      -- CP-element group 342: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/type_cast_1115_Sample/ra
      -- 
    ra_2638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 342_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1115_inst_ack_0, ack => convTranspose_CP_39_elements(342)); -- 
    -- CP-element group 343:  transition  input  output  bypass 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	339 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	344 
    -- CP-element group 343:  members (6) 
      -- CP-element group 343: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/type_cast_1115_update_completed_
      -- CP-element group 343: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/type_cast_1115_Update/$exit
      -- CP-element group 343: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/type_cast_1115_Update/ca
      -- CP-element group 343: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/WPIPE_elapsed_time_pipe_1122_sample_start_
      -- CP-element group 343: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/WPIPE_elapsed_time_pipe_1122_Sample/$entry
      -- CP-element group 343: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/WPIPE_elapsed_time_pipe_1122_Sample/req
      -- 
    ca_2643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 343_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1115_inst_ack_1, ack => convTranspose_CP_39_elements(343)); -- 
    req_2651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(343), ack => WPIPE_elapsed_time_pipe_1122_inst_req_0); -- 
    -- CP-element group 344:  transition  input  output  bypass 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	343 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	345 
    -- CP-element group 344:  members (6) 
      -- CP-element group 344: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/WPIPE_elapsed_time_pipe_1122_sample_completed_
      -- CP-element group 344: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/WPIPE_elapsed_time_pipe_1122_update_start_
      -- CP-element group 344: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/WPIPE_elapsed_time_pipe_1122_Sample/$exit
      -- CP-element group 344: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/WPIPE_elapsed_time_pipe_1122_Sample/ack
      -- CP-element group 344: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/WPIPE_elapsed_time_pipe_1122_Update/$entry
      -- CP-element group 344: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/WPIPE_elapsed_time_pipe_1122_Update/req
      -- 
    ack_2652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 344_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1122_inst_ack_0, ack => convTranspose_CP_39_elements(344)); -- 
    req_2656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(344), ack => WPIPE_elapsed_time_pipe_1122_inst_req_1); -- 
    -- CP-element group 345:  branch  transition  place  input  output  bypass 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	344 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	346 
    -- CP-element group 345: 	347 
    -- CP-element group 345:  members (13) 
      -- CP-element group 345: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124__exit__
      -- CP-element group 345: 	 branch_block_stmt_33/if_stmt_1126__entry__
      -- CP-element group 345: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/$exit
      -- CP-element group 345: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/WPIPE_elapsed_time_pipe_1122_update_completed_
      -- CP-element group 345: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/WPIPE_elapsed_time_pipe_1122_Update/$exit
      -- CP-element group 345: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/WPIPE_elapsed_time_pipe_1122_Update/ack
      -- CP-element group 345: 	 branch_block_stmt_33/if_stmt_1126_dead_link/$entry
      -- CP-element group 345: 	 branch_block_stmt_33/if_stmt_1126_eval_test/$entry
      -- CP-element group 345: 	 branch_block_stmt_33/if_stmt_1126_eval_test/$exit
      -- CP-element group 345: 	 branch_block_stmt_33/if_stmt_1126_eval_test/branch_req
      -- CP-element group 345: 	 branch_block_stmt_33/R_cmp250409_1127_place
      -- CP-element group 345: 	 branch_block_stmt_33/if_stmt_1126_if_link/$entry
      -- CP-element group 345: 	 branch_block_stmt_33/if_stmt_1126_else_link/$entry
      -- 
    ack_2657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 345_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1122_inst_ack_1, ack => convTranspose_CP_39_elements(345)); -- 
    branch_req_2665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(345), ack => if_stmt_1126_branch_req_0); -- 
    -- CP-element group 346:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	345 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	348 
    -- CP-element group 346: 	349 
    -- CP-element group 346:  members (18) 
      -- CP-element group 346: 	 branch_block_stmt_33/merge_stmt_1132__exit__
      -- CP-element group 346: 	 branch_block_stmt_33/assign_stmt_1138_to_assign_stmt_1167__entry__
      -- CP-element group 346: 	 branch_block_stmt_33/merge_stmt_1132_PhiAck/dummy
      -- CP-element group 346: 	 branch_block_stmt_33/merge_stmt_1132_PhiAck/$exit
      -- CP-element group 346: 	 branch_block_stmt_33/merge_stmt_1132_PhiReqMerge
      -- CP-element group 346: 	 branch_block_stmt_33/merge_stmt_1132_PhiAck/$entry
      -- CP-element group 346: 	 branch_block_stmt_33/forx_xend259_bbx_xnph_PhiReq/$exit
      -- CP-element group 346: 	 branch_block_stmt_33/forx_xend259_bbx_xnph_PhiReq/$entry
      -- CP-element group 346: 	 branch_block_stmt_33/if_stmt_1126_if_link/$exit
      -- CP-element group 346: 	 branch_block_stmt_33/if_stmt_1126_if_link/if_choice_transition
      -- CP-element group 346: 	 branch_block_stmt_33/forx_xend259_bbx_xnph
      -- CP-element group 346: 	 branch_block_stmt_33/assign_stmt_1138_to_assign_stmt_1167/$entry
      -- CP-element group 346: 	 branch_block_stmt_33/assign_stmt_1138_to_assign_stmt_1167/type_cast_1153_sample_start_
      -- CP-element group 346: 	 branch_block_stmt_33/assign_stmt_1138_to_assign_stmt_1167/type_cast_1153_update_start_
      -- CP-element group 346: 	 branch_block_stmt_33/assign_stmt_1138_to_assign_stmt_1167/type_cast_1153_Sample/$entry
      -- CP-element group 346: 	 branch_block_stmt_33/assign_stmt_1138_to_assign_stmt_1167/type_cast_1153_Sample/rr
      -- CP-element group 346: 	 branch_block_stmt_33/assign_stmt_1138_to_assign_stmt_1167/type_cast_1153_Update/$entry
      -- CP-element group 346: 	 branch_block_stmt_33/assign_stmt_1138_to_assign_stmt_1167/type_cast_1153_Update/cr
      -- 
    if_choice_transition_2670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 346_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1126_branch_ack_1, ack => convTranspose_CP_39_elements(346)); -- 
    rr_2687_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2687_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(346), ack => type_cast_1153_inst_req_0); -- 
    cr_2692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(346), ack => type_cast_1153_inst_req_1); -- 
    -- CP-element group 347:  transition  place  input  bypass 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	345 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	425 
    -- CP-element group 347:  members (5) 
      -- CP-element group 347: 	 branch_block_stmt_33/forx_xend259_forx_xend404_PhiReq/$exit
      -- CP-element group 347: 	 branch_block_stmt_33/forx_xend259_forx_xend404_PhiReq/$entry
      -- CP-element group 347: 	 branch_block_stmt_33/if_stmt_1126_else_link/$exit
      -- CP-element group 347: 	 branch_block_stmt_33/if_stmt_1126_else_link/else_choice_transition
      -- CP-element group 347: 	 branch_block_stmt_33/forx_xend259_forx_xend404
      -- 
    else_choice_transition_2674_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 347_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1126_branch_ack_0, ack => convTranspose_CP_39_elements(347)); -- 
    -- CP-element group 348:  transition  input  bypass 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	346 
    -- CP-element group 348: successors 
    -- CP-element group 348:  members (3) 
      -- CP-element group 348: 	 branch_block_stmt_33/assign_stmt_1138_to_assign_stmt_1167/type_cast_1153_sample_completed_
      -- CP-element group 348: 	 branch_block_stmt_33/assign_stmt_1138_to_assign_stmt_1167/type_cast_1153_Sample/$exit
      -- CP-element group 348: 	 branch_block_stmt_33/assign_stmt_1138_to_assign_stmt_1167/type_cast_1153_Sample/ra
      -- 
    ra_2688_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 348_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1153_inst_ack_0, ack => convTranspose_CP_39_elements(348)); -- 
    -- CP-element group 349:  transition  place  input  bypass 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	346 
    -- CP-element group 349: successors 
    -- CP-element group 349: 	419 
    -- CP-element group 349:  members (9) 
      -- CP-element group 349: 	 branch_block_stmt_33/assign_stmt_1138_to_assign_stmt_1167__exit__
      -- CP-element group 349: 	 branch_block_stmt_33/bbx_xnph_forx_xbody332
      -- CP-element group 349: 	 branch_block_stmt_33/bbx_xnph_forx_xbody332_PhiReq/$entry
      -- CP-element group 349: 	 branch_block_stmt_33/bbx_xnph_forx_xbody332_PhiReq/phi_stmt_1170/$entry
      -- CP-element group 349: 	 branch_block_stmt_33/bbx_xnph_forx_xbody332_PhiReq/phi_stmt_1170/phi_stmt_1170_sources/$entry
      -- CP-element group 349: 	 branch_block_stmt_33/assign_stmt_1138_to_assign_stmt_1167/$exit
      -- CP-element group 349: 	 branch_block_stmt_33/assign_stmt_1138_to_assign_stmt_1167/type_cast_1153_update_completed_
      -- CP-element group 349: 	 branch_block_stmt_33/assign_stmt_1138_to_assign_stmt_1167/type_cast_1153_Update/$exit
      -- CP-element group 349: 	 branch_block_stmt_33/assign_stmt_1138_to_assign_stmt_1167/type_cast_1153_Update/ca
      -- 
    ca_2693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 349_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1153_inst_ack_1, ack => convTranspose_CP_39_elements(349)); -- 
    -- CP-element group 350:  transition  input  bypass 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	424 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	395 
    -- CP-element group 350:  members (3) 
      -- CP-element group 350: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/array_obj_ref_1182_final_index_sum_regn_sample_complete
      -- CP-element group 350: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/array_obj_ref_1182_final_index_sum_regn_Sample/$exit
      -- CP-element group 350: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/array_obj_ref_1182_final_index_sum_regn_Sample/ack
      -- 
    ack_2722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 350_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1182_index_offset_ack_0, ack => convTranspose_CP_39_elements(350)); -- 
    -- CP-element group 351:  transition  input  output  bypass 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	424 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	352 
    -- CP-element group 351:  members (11) 
      -- CP-element group 351: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/addr_of_1183_sample_start_
      -- CP-element group 351: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/array_obj_ref_1182_root_address_calculated
      -- CP-element group 351: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/array_obj_ref_1182_offset_calculated
      -- CP-element group 351: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/array_obj_ref_1182_final_index_sum_regn_Update/$exit
      -- CP-element group 351: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/array_obj_ref_1182_final_index_sum_regn_Update/ack
      -- CP-element group 351: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/array_obj_ref_1182_base_plus_offset/$entry
      -- CP-element group 351: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/array_obj_ref_1182_base_plus_offset/$exit
      -- CP-element group 351: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/array_obj_ref_1182_base_plus_offset/sum_rename_req
      -- CP-element group 351: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/array_obj_ref_1182_base_plus_offset/sum_rename_ack
      -- CP-element group 351: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/addr_of_1183_request/$entry
      -- CP-element group 351: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/addr_of_1183_request/req
      -- 
    ack_2727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 351_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1182_index_offset_ack_1, ack => convTranspose_CP_39_elements(351)); -- 
    req_2736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(351), ack => addr_of_1183_final_reg_req_0); -- 
    -- CP-element group 352:  transition  input  bypass 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	351 
    -- CP-element group 352: successors 
    -- CP-element group 352:  members (3) 
      -- CP-element group 352: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/addr_of_1183_sample_completed_
      -- CP-element group 352: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/addr_of_1183_request/$exit
      -- CP-element group 352: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/addr_of_1183_request/ack
      -- 
    ack_2737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1183_final_reg_ack_0, ack => convTranspose_CP_39_elements(352)); -- 
    -- CP-element group 353:  join  fork  transition  input  output  bypass 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	424 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	354 
    -- CP-element group 353:  members (24) 
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/addr_of_1183_update_completed_
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/addr_of_1183_complete/$exit
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/addr_of_1183_complete/ack
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/ptr_deref_1187_sample_start_
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/ptr_deref_1187_base_address_calculated
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/ptr_deref_1187_word_address_calculated
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/ptr_deref_1187_root_address_calculated
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/ptr_deref_1187_base_address_resized
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/ptr_deref_1187_base_addr_resize/$entry
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/ptr_deref_1187_base_addr_resize/$exit
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/ptr_deref_1187_base_addr_resize/base_resize_req
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/ptr_deref_1187_base_addr_resize/base_resize_ack
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/ptr_deref_1187_base_plus_offset/$entry
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/ptr_deref_1187_base_plus_offset/$exit
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/ptr_deref_1187_base_plus_offset/sum_rename_req
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/ptr_deref_1187_base_plus_offset/sum_rename_ack
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/ptr_deref_1187_word_addrgen/$entry
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/ptr_deref_1187_word_addrgen/$exit
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/ptr_deref_1187_word_addrgen/root_register_req
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/ptr_deref_1187_word_addrgen/root_register_ack
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/ptr_deref_1187_Sample/$entry
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/ptr_deref_1187_Sample/word_access_start/$entry
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/ptr_deref_1187_Sample/word_access_start/word_0/$entry
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/ptr_deref_1187_Sample/word_access_start/word_0/rr
      -- 
    ack_2742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 353_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1183_final_reg_ack_1, ack => convTranspose_CP_39_elements(353)); -- 
    rr_2775_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2775_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(353), ack => ptr_deref_1187_load_0_req_0); -- 
    -- CP-element group 354:  transition  input  bypass 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	353 
    -- CP-element group 354: successors 
    -- CP-element group 354:  members (5) 
      -- CP-element group 354: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/ptr_deref_1187_sample_completed_
      -- CP-element group 354: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/ptr_deref_1187_Sample/$exit
      -- CP-element group 354: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/ptr_deref_1187_Sample/word_access_start/$exit
      -- CP-element group 354: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/ptr_deref_1187_Sample/word_access_start/word_0/$exit
      -- CP-element group 354: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/ptr_deref_1187_Sample/word_access_start/word_0/ra
      -- 
    ra_2776_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 354_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1187_load_0_ack_0, ack => convTranspose_CP_39_elements(354)); -- 
    -- CP-element group 355:  fork  transition  input  output  bypass 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	424 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	356 
    -- CP-element group 355: 	358 
    -- CP-element group 355: 	360 
    -- CP-element group 355: 	362 
    -- CP-element group 355: 	364 
    -- CP-element group 355: 	366 
    -- CP-element group 355: 	368 
    -- CP-element group 355: 	370 
    -- CP-element group 355:  members (33) 
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/ptr_deref_1187_update_completed_
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/ptr_deref_1187_Update/$exit
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/ptr_deref_1187_Update/word_access_complete/$exit
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/ptr_deref_1187_Update/word_access_complete/word_0/$exit
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/ptr_deref_1187_Update/word_access_complete/word_0/ca
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/ptr_deref_1187_Update/ptr_deref_1187_Merge/$entry
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/ptr_deref_1187_Update/ptr_deref_1187_Merge/$exit
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/ptr_deref_1187_Update/ptr_deref_1187_Merge/merge_req
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/ptr_deref_1187_Update/ptr_deref_1187_Merge/merge_ack
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1191_sample_start_
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1191_Sample/$entry
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1191_Sample/rr
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1201_sample_start_
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1201_Sample/$entry
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1201_Sample/rr
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1211_sample_start_
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1211_Sample/$entry
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1211_Sample/rr
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1221_sample_start_
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1221_Sample/$entry
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1221_Sample/rr
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1231_sample_start_
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1231_Sample/$entry
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1231_Sample/rr
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1241_sample_start_
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1241_Sample/$entry
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1241_Sample/rr
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1251_sample_start_
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1251_Sample/$entry
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1251_Sample/rr
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1261_sample_start_
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1261_Sample/$entry
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1261_Sample/rr
      -- 
    ca_2787_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 355_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1187_load_0_ack_1, ack => convTranspose_CP_39_elements(355)); -- 
    rr_2800_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2800_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(355), ack => type_cast_1191_inst_req_0); -- 
    rr_2814_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2814_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(355), ack => type_cast_1201_inst_req_0); -- 
    rr_2828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(355), ack => type_cast_1211_inst_req_0); -- 
    rr_2842_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2842_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(355), ack => type_cast_1221_inst_req_0); -- 
    rr_2856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(355), ack => type_cast_1231_inst_req_0); -- 
    rr_2870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(355), ack => type_cast_1241_inst_req_0); -- 
    rr_2884_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2884_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(355), ack => type_cast_1251_inst_req_0); -- 
    rr_2898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(355), ack => type_cast_1261_inst_req_0); -- 
    -- CP-element group 356:  transition  input  bypass 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	355 
    -- CP-element group 356: successors 
    -- CP-element group 356:  members (3) 
      -- CP-element group 356: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1191_sample_completed_
      -- CP-element group 356: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1191_Sample/$exit
      -- CP-element group 356: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1191_Sample/ra
      -- 
    ra_2801_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 356_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1191_inst_ack_0, ack => convTranspose_CP_39_elements(356)); -- 
    -- CP-element group 357:  transition  input  bypass 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	424 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	392 
    -- CP-element group 357:  members (3) 
      -- CP-element group 357: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1191_update_completed_
      -- CP-element group 357: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1191_Update/$exit
      -- CP-element group 357: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1191_Update/ca
      -- 
    ca_2806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 357_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1191_inst_ack_1, ack => convTranspose_CP_39_elements(357)); -- 
    -- CP-element group 358:  transition  input  bypass 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	355 
    -- CP-element group 358: successors 
    -- CP-element group 358:  members (3) 
      -- CP-element group 358: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1201_sample_completed_
      -- CP-element group 358: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1201_Sample/$exit
      -- CP-element group 358: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1201_Sample/ra
      -- 
    ra_2815_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 358_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1201_inst_ack_0, ack => convTranspose_CP_39_elements(358)); -- 
    -- CP-element group 359:  transition  input  bypass 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	424 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	389 
    -- CP-element group 359:  members (3) 
      -- CP-element group 359: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1201_update_completed_
      -- CP-element group 359: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1201_Update/$exit
      -- CP-element group 359: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1201_Update/ca
      -- 
    ca_2820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 359_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1201_inst_ack_1, ack => convTranspose_CP_39_elements(359)); -- 
    -- CP-element group 360:  transition  input  bypass 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	355 
    -- CP-element group 360: successors 
    -- CP-element group 360:  members (3) 
      -- CP-element group 360: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1211_sample_completed_
      -- CP-element group 360: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1211_Sample/$exit
      -- CP-element group 360: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1211_Sample/ra
      -- 
    ra_2829_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 360_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1211_inst_ack_0, ack => convTranspose_CP_39_elements(360)); -- 
    -- CP-element group 361:  transition  input  bypass 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	424 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	386 
    -- CP-element group 361:  members (3) 
      -- CP-element group 361: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1211_update_completed_
      -- CP-element group 361: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1211_Update/$exit
      -- CP-element group 361: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1211_Update/ca
      -- 
    ca_2834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 361_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1211_inst_ack_1, ack => convTranspose_CP_39_elements(361)); -- 
    -- CP-element group 362:  transition  input  bypass 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	355 
    -- CP-element group 362: successors 
    -- CP-element group 362:  members (3) 
      -- CP-element group 362: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1221_sample_completed_
      -- CP-element group 362: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1221_Sample/$exit
      -- CP-element group 362: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1221_Sample/ra
      -- 
    ra_2843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 362_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1221_inst_ack_0, ack => convTranspose_CP_39_elements(362)); -- 
    -- CP-element group 363:  transition  input  bypass 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	424 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	383 
    -- CP-element group 363:  members (3) 
      -- CP-element group 363: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1221_update_completed_
      -- CP-element group 363: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1221_Update/$exit
      -- CP-element group 363: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1221_Update/ca
      -- 
    ca_2848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 363_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1221_inst_ack_1, ack => convTranspose_CP_39_elements(363)); -- 
    -- CP-element group 364:  transition  input  bypass 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	355 
    -- CP-element group 364: successors 
    -- CP-element group 364:  members (3) 
      -- CP-element group 364: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1231_sample_completed_
      -- CP-element group 364: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1231_Sample/$exit
      -- CP-element group 364: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1231_Sample/ra
      -- 
    ra_2857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 364_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1231_inst_ack_0, ack => convTranspose_CP_39_elements(364)); -- 
    -- CP-element group 365:  transition  input  bypass 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	424 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	380 
    -- CP-element group 365:  members (3) 
      -- CP-element group 365: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1231_update_completed_
      -- CP-element group 365: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1231_Update/$exit
      -- CP-element group 365: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1231_Update/ca
      -- 
    ca_2862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 365_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1231_inst_ack_1, ack => convTranspose_CP_39_elements(365)); -- 
    -- CP-element group 366:  transition  input  bypass 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	355 
    -- CP-element group 366: successors 
    -- CP-element group 366:  members (3) 
      -- CP-element group 366: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1241_sample_completed_
      -- CP-element group 366: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1241_Sample/$exit
      -- CP-element group 366: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1241_Sample/ra
      -- 
    ra_2871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 366_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1241_inst_ack_0, ack => convTranspose_CP_39_elements(366)); -- 
    -- CP-element group 367:  transition  input  bypass 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	424 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	377 
    -- CP-element group 367:  members (3) 
      -- CP-element group 367: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1241_update_completed_
      -- CP-element group 367: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1241_Update/$exit
      -- CP-element group 367: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1241_Update/ca
      -- 
    ca_2876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 367_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1241_inst_ack_1, ack => convTranspose_CP_39_elements(367)); -- 
    -- CP-element group 368:  transition  input  bypass 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	355 
    -- CP-element group 368: successors 
    -- CP-element group 368:  members (3) 
      -- CP-element group 368: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1251_sample_completed_
      -- CP-element group 368: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1251_Sample/$exit
      -- CP-element group 368: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1251_Sample/ra
      -- 
    ra_2885_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 368_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1251_inst_ack_0, ack => convTranspose_CP_39_elements(368)); -- 
    -- CP-element group 369:  transition  input  bypass 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	424 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	374 
    -- CP-element group 369:  members (3) 
      -- CP-element group 369: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1251_update_completed_
      -- CP-element group 369: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1251_Update/$exit
      -- CP-element group 369: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1251_Update/ca
      -- 
    ca_2890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 369_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1251_inst_ack_1, ack => convTranspose_CP_39_elements(369)); -- 
    -- CP-element group 370:  transition  input  bypass 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	355 
    -- CP-element group 370: successors 
    -- CP-element group 370:  members (3) 
      -- CP-element group 370: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1261_sample_completed_
      -- CP-element group 370: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1261_Sample/$exit
      -- CP-element group 370: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1261_Sample/ra
      -- 
    ra_2899_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 370_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1261_inst_ack_0, ack => convTranspose_CP_39_elements(370)); -- 
    -- CP-element group 371:  transition  input  output  bypass 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	424 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	372 
    -- CP-element group 371:  members (6) 
      -- CP-element group 371: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1261_update_completed_
      -- CP-element group 371: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1261_Update/$exit
      -- CP-element group 371: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1261_Update/ca
      -- CP-element group 371: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1263_sample_start_
      -- CP-element group 371: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1263_Sample/$entry
      -- CP-element group 371: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1263_Sample/req
      -- 
    ca_2904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 371_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1261_inst_ack_1, ack => convTranspose_CP_39_elements(371)); -- 
    req_2912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(371), ack => WPIPE_ConvTranspose_output_pipe_1263_inst_req_0); -- 
    -- CP-element group 372:  transition  input  output  bypass 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	371 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	373 
    -- CP-element group 372:  members (6) 
      -- CP-element group 372: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1263_sample_completed_
      -- CP-element group 372: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1263_update_start_
      -- CP-element group 372: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1263_Sample/$exit
      -- CP-element group 372: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1263_Sample/ack
      -- CP-element group 372: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1263_Update/$entry
      -- CP-element group 372: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1263_Update/req
      -- 
    ack_2913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 372_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1263_inst_ack_0, ack => convTranspose_CP_39_elements(372)); -- 
    req_2917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(372), ack => WPIPE_ConvTranspose_output_pipe_1263_inst_req_1); -- 
    -- CP-element group 373:  transition  input  bypass 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	372 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	374 
    -- CP-element group 373:  members (3) 
      -- CP-element group 373: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1263_update_completed_
      -- CP-element group 373: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1263_Update/$exit
      -- CP-element group 373: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1263_Update/ack
      -- 
    ack_2918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 373_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1263_inst_ack_1, ack => convTranspose_CP_39_elements(373)); -- 
    -- CP-element group 374:  join  transition  output  bypass 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	369 
    -- CP-element group 374: 	373 
    -- CP-element group 374: successors 
    -- CP-element group 374: 	375 
    -- CP-element group 374:  members (3) 
      -- CP-element group 374: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1266_sample_start_
      -- CP-element group 374: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1266_Sample/$entry
      -- CP-element group 374: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1266_Sample/req
      -- 
    req_2926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(374), ack => WPIPE_ConvTranspose_output_pipe_1266_inst_req_0); -- 
    convTranspose_cp_element_group_374: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_374"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(369) & convTranspose_CP_39_elements(373);
      gj_convTranspose_cp_element_group_374 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(374), clk => clk, reset => reset); --
    end block;
    -- CP-element group 375:  transition  input  output  bypass 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	374 
    -- CP-element group 375: successors 
    -- CP-element group 375: 	376 
    -- CP-element group 375:  members (6) 
      -- CP-element group 375: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1266_sample_completed_
      -- CP-element group 375: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1266_update_start_
      -- CP-element group 375: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1266_Sample/$exit
      -- CP-element group 375: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1266_Sample/ack
      -- CP-element group 375: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1266_Update/$entry
      -- CP-element group 375: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1266_Update/req
      -- 
    ack_2927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 375_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1266_inst_ack_0, ack => convTranspose_CP_39_elements(375)); -- 
    req_2931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(375), ack => WPIPE_ConvTranspose_output_pipe_1266_inst_req_1); -- 
    -- CP-element group 376:  transition  input  bypass 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	375 
    -- CP-element group 376: successors 
    -- CP-element group 376: 	377 
    -- CP-element group 376:  members (3) 
      -- CP-element group 376: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1266_update_completed_
      -- CP-element group 376: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1266_Update/$exit
      -- CP-element group 376: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1266_Update/ack
      -- 
    ack_2932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 376_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1266_inst_ack_1, ack => convTranspose_CP_39_elements(376)); -- 
    -- CP-element group 377:  join  transition  output  bypass 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	367 
    -- CP-element group 377: 	376 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	378 
    -- CP-element group 377:  members (3) 
      -- CP-element group 377: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1269_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1269_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1269_Sample/req
      -- 
    req_2940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(377), ack => WPIPE_ConvTranspose_output_pipe_1269_inst_req_0); -- 
    convTranspose_cp_element_group_377: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_377"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(367) & convTranspose_CP_39_elements(376);
      gj_convTranspose_cp_element_group_377 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(377), clk => clk, reset => reset); --
    end block;
    -- CP-element group 378:  transition  input  output  bypass 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	377 
    -- CP-element group 378: successors 
    -- CP-element group 378: 	379 
    -- CP-element group 378:  members (6) 
      -- CP-element group 378: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1269_sample_completed_
      -- CP-element group 378: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1269_update_start_
      -- CP-element group 378: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1269_Sample/$exit
      -- CP-element group 378: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1269_Sample/ack
      -- CP-element group 378: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1269_Update/$entry
      -- CP-element group 378: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1269_Update/req
      -- 
    ack_2941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 378_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1269_inst_ack_0, ack => convTranspose_CP_39_elements(378)); -- 
    req_2945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(378), ack => WPIPE_ConvTranspose_output_pipe_1269_inst_req_1); -- 
    -- CP-element group 379:  transition  input  bypass 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	378 
    -- CP-element group 379: successors 
    -- CP-element group 379: 	380 
    -- CP-element group 379:  members (3) 
      -- CP-element group 379: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1269_update_completed_
      -- CP-element group 379: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1269_Update/$exit
      -- CP-element group 379: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1269_Update/ack
      -- 
    ack_2946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 379_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1269_inst_ack_1, ack => convTranspose_CP_39_elements(379)); -- 
    -- CP-element group 380:  join  transition  output  bypass 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	365 
    -- CP-element group 380: 	379 
    -- CP-element group 380: successors 
    -- CP-element group 380: 	381 
    -- CP-element group 380:  members (3) 
      -- CP-element group 380: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1272_sample_start_
      -- CP-element group 380: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1272_Sample/$entry
      -- CP-element group 380: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1272_Sample/req
      -- 
    req_2954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(380), ack => WPIPE_ConvTranspose_output_pipe_1272_inst_req_0); -- 
    convTranspose_cp_element_group_380: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_380"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(365) & convTranspose_CP_39_elements(379);
      gj_convTranspose_cp_element_group_380 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(380), clk => clk, reset => reset); --
    end block;
    -- CP-element group 381:  transition  input  output  bypass 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	380 
    -- CP-element group 381: successors 
    -- CP-element group 381: 	382 
    -- CP-element group 381:  members (6) 
      -- CP-element group 381: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1272_sample_completed_
      -- CP-element group 381: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1272_update_start_
      -- CP-element group 381: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1272_Sample/$exit
      -- CP-element group 381: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1272_Sample/ack
      -- CP-element group 381: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1272_Update/$entry
      -- CP-element group 381: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1272_Update/req
      -- 
    ack_2955_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 381_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1272_inst_ack_0, ack => convTranspose_CP_39_elements(381)); -- 
    req_2959_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2959_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(381), ack => WPIPE_ConvTranspose_output_pipe_1272_inst_req_1); -- 
    -- CP-element group 382:  transition  input  bypass 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	381 
    -- CP-element group 382: successors 
    -- CP-element group 382: 	383 
    -- CP-element group 382:  members (3) 
      -- CP-element group 382: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1272_update_completed_
      -- CP-element group 382: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1272_Update/$exit
      -- CP-element group 382: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1272_Update/ack
      -- 
    ack_2960_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 382_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1272_inst_ack_1, ack => convTranspose_CP_39_elements(382)); -- 
    -- CP-element group 383:  join  transition  output  bypass 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	363 
    -- CP-element group 383: 	382 
    -- CP-element group 383: successors 
    -- CP-element group 383: 	384 
    -- CP-element group 383:  members (3) 
      -- CP-element group 383: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1275_sample_start_
      -- CP-element group 383: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1275_Sample/$entry
      -- CP-element group 383: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1275_Sample/req
      -- 
    req_2968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(383), ack => WPIPE_ConvTranspose_output_pipe_1275_inst_req_0); -- 
    convTranspose_cp_element_group_383: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_383"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(363) & convTranspose_CP_39_elements(382);
      gj_convTranspose_cp_element_group_383 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(383), clk => clk, reset => reset); --
    end block;
    -- CP-element group 384:  transition  input  output  bypass 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	383 
    -- CP-element group 384: successors 
    -- CP-element group 384: 	385 
    -- CP-element group 384:  members (6) 
      -- CP-element group 384: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1275_Update/req
      -- CP-element group 384: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1275_sample_completed_
      -- CP-element group 384: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1275_update_start_
      -- CP-element group 384: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1275_Sample/$exit
      -- CP-element group 384: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1275_Sample/ack
      -- CP-element group 384: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1275_Update/$entry
      -- 
    ack_2969_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 384_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1275_inst_ack_0, ack => convTranspose_CP_39_elements(384)); -- 
    req_2973_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2973_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(384), ack => WPIPE_ConvTranspose_output_pipe_1275_inst_req_1); -- 
    -- CP-element group 385:  transition  input  bypass 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	384 
    -- CP-element group 385: successors 
    -- CP-element group 385: 	386 
    -- CP-element group 385:  members (3) 
      -- CP-element group 385: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1275_Update/ack
      -- CP-element group 385: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1275_Update/$exit
      -- CP-element group 385: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1275_update_completed_
      -- 
    ack_2974_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 385_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1275_inst_ack_1, ack => convTranspose_CP_39_elements(385)); -- 
    -- CP-element group 386:  join  transition  output  bypass 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	361 
    -- CP-element group 386: 	385 
    -- CP-element group 386: successors 
    -- CP-element group 386: 	387 
    -- CP-element group 386:  members (3) 
      -- CP-element group 386: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1278_sample_start_
      -- CP-element group 386: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1278_Sample/$entry
      -- CP-element group 386: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1278_Sample/req
      -- 
    req_2982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(386), ack => WPIPE_ConvTranspose_output_pipe_1278_inst_req_0); -- 
    convTranspose_cp_element_group_386: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_386"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(361) & convTranspose_CP_39_elements(385);
      gj_convTranspose_cp_element_group_386 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(386), clk => clk, reset => reset); --
    end block;
    -- CP-element group 387:  transition  input  output  bypass 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	386 
    -- CP-element group 387: successors 
    -- CP-element group 387: 	388 
    -- CP-element group 387:  members (6) 
      -- CP-element group 387: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1278_sample_completed_
      -- CP-element group 387: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1278_update_start_
      -- CP-element group 387: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1278_Sample/$exit
      -- CP-element group 387: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1278_Sample/ack
      -- CP-element group 387: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1278_Update/$entry
      -- CP-element group 387: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1278_Update/req
      -- 
    ack_2983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 387_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1278_inst_ack_0, ack => convTranspose_CP_39_elements(387)); -- 
    req_2987_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2987_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(387), ack => WPIPE_ConvTranspose_output_pipe_1278_inst_req_1); -- 
    -- CP-element group 388:  transition  input  bypass 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: 	387 
    -- CP-element group 388: successors 
    -- CP-element group 388: 	389 
    -- CP-element group 388:  members (3) 
      -- CP-element group 388: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1278_update_completed_
      -- CP-element group 388: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1278_Update/$exit
      -- CP-element group 388: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1278_Update/ack
      -- 
    ack_2988_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 388_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1278_inst_ack_1, ack => convTranspose_CP_39_elements(388)); -- 
    -- CP-element group 389:  join  transition  output  bypass 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	359 
    -- CP-element group 389: 	388 
    -- CP-element group 389: successors 
    -- CP-element group 389: 	390 
    -- CP-element group 389:  members (3) 
      -- CP-element group 389: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1281_Sample/req
      -- CP-element group 389: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1281_Sample/$entry
      -- CP-element group 389: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1281_sample_start_
      -- 
    req_2996_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2996_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(389), ack => WPIPE_ConvTranspose_output_pipe_1281_inst_req_0); -- 
    convTranspose_cp_element_group_389: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_389"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(359) & convTranspose_CP_39_elements(388);
      gj_convTranspose_cp_element_group_389 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(389), clk => clk, reset => reset); --
    end block;
    -- CP-element group 390:  transition  input  output  bypass 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: 	389 
    -- CP-element group 390: successors 
    -- CP-element group 390: 	391 
    -- CP-element group 390:  members (6) 
      -- CP-element group 390: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1281_Sample/ack
      -- CP-element group 390: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1281_Update/$entry
      -- CP-element group 390: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1281_Update/req
      -- CP-element group 390: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1281_Sample/$exit
      -- CP-element group 390: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1281_update_start_
      -- CP-element group 390: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1281_sample_completed_
      -- 
    ack_2997_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 390_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1281_inst_ack_0, ack => convTranspose_CP_39_elements(390)); -- 
    req_3001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(390), ack => WPIPE_ConvTranspose_output_pipe_1281_inst_req_1); -- 
    -- CP-element group 391:  transition  input  bypass 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: 	390 
    -- CP-element group 391: successors 
    -- CP-element group 391: 	392 
    -- CP-element group 391:  members (3) 
      -- CP-element group 391: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1281_Update/$exit
      -- CP-element group 391: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1281_Update/ack
      -- CP-element group 391: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1281_update_completed_
      -- 
    ack_3002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 391_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1281_inst_ack_1, ack => convTranspose_CP_39_elements(391)); -- 
    -- CP-element group 392:  join  transition  output  bypass 
    -- CP-element group 392: predecessors 
    -- CP-element group 392: 	357 
    -- CP-element group 392: 	391 
    -- CP-element group 392: successors 
    -- CP-element group 392: 	393 
    -- CP-element group 392:  members (3) 
      -- CP-element group 392: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1284_sample_start_
      -- CP-element group 392: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1284_Sample/req
      -- CP-element group 392: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1284_Sample/$entry
      -- 
    req_3010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(392), ack => WPIPE_ConvTranspose_output_pipe_1284_inst_req_0); -- 
    convTranspose_cp_element_group_392: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_392"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(357) & convTranspose_CP_39_elements(391);
      gj_convTranspose_cp_element_group_392 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(392), clk => clk, reset => reset); --
    end block;
    -- CP-element group 393:  transition  input  output  bypass 
    -- CP-element group 393: predecessors 
    -- CP-element group 393: 	392 
    -- CP-element group 393: successors 
    -- CP-element group 393: 	394 
    -- CP-element group 393:  members (6) 
      -- CP-element group 393: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1284_sample_completed_
      -- CP-element group 393: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1284_Update/req
      -- CP-element group 393: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1284_Update/$entry
      -- CP-element group 393: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1284_Sample/ack
      -- CP-element group 393: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1284_Sample/$exit
      -- CP-element group 393: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1284_update_start_
      -- 
    ack_3011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 393_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1284_inst_ack_0, ack => convTranspose_CP_39_elements(393)); -- 
    req_3015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(393), ack => WPIPE_ConvTranspose_output_pipe_1284_inst_req_1); -- 
    -- CP-element group 394:  transition  input  bypass 
    -- CP-element group 394: predecessors 
    -- CP-element group 394: 	393 
    -- CP-element group 394: successors 
    -- CP-element group 394: 	395 
    -- CP-element group 394:  members (3) 
      -- CP-element group 394: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1284_Update/ack
      -- CP-element group 394: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1284_Update/$exit
      -- CP-element group 394: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/WPIPE_ConvTranspose_output_pipe_1284_update_completed_
      -- 
    ack_3016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 394_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1284_inst_ack_1, ack => convTranspose_CP_39_elements(394)); -- 
    -- CP-element group 395:  branch  join  transition  place  output  bypass 
    -- CP-element group 395: predecessors 
    -- CP-element group 395: 	350 
    -- CP-element group 395: 	394 
    -- CP-element group 395: successors 
    -- CP-element group 395: 	396 
    -- CP-element group 395: 	397 
    -- CP-element group 395:  members (10) 
      -- CP-element group 395: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297__exit__
      -- CP-element group 395: 	 branch_block_stmt_33/if_stmt_1298__entry__
      -- CP-element group 395: 	 branch_block_stmt_33/if_stmt_1298_else_link/$entry
      -- CP-element group 395: 	 branch_block_stmt_33/if_stmt_1298_if_link/$entry
      -- CP-element group 395: 	 branch_block_stmt_33/if_stmt_1298_eval_test/$exit
      -- CP-element group 395: 	 branch_block_stmt_33/if_stmt_1298_eval_test/branch_req
      -- CP-element group 395: 	 branch_block_stmt_33/if_stmt_1298_eval_test/$entry
      -- CP-element group 395: 	 branch_block_stmt_33/if_stmt_1298_dead_link/$entry
      -- CP-element group 395: 	 branch_block_stmt_33/R_exitcond1_1299_place
      -- CP-element group 395: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/$exit
      -- 
    branch_req_3024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(395), ack => if_stmt_1298_branch_req_0); -- 
    convTranspose_cp_element_group_395: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_395"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(350) & convTranspose_CP_39_elements(394);
      gj_convTranspose_cp_element_group_395 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(395), clk => clk, reset => reset); --
    end block;
    -- CP-element group 396:  merge  transition  place  input  bypass 
    -- CP-element group 396: predecessors 
    -- CP-element group 396: 	395 
    -- CP-element group 396: successors 
    -- CP-element group 396: 	425 
    -- CP-element group 396:  members (13) 
      -- CP-element group 396: 	 branch_block_stmt_33/if_stmt_1298_if_link/$exit
      -- CP-element group 396: 	 branch_block_stmt_33/merge_stmt_1304__exit__
      -- CP-element group 396: 	 branch_block_stmt_33/forx_xend404x_xloopexit_forx_xend404
      -- CP-element group 396: 	 branch_block_stmt_33/if_stmt_1298_if_link/if_choice_transition
      -- CP-element group 396: 	 branch_block_stmt_33/forx_xend404x_xloopexit_forx_xend404_PhiReq/$exit
      -- CP-element group 396: 	 branch_block_stmt_33/merge_stmt_1304_PhiReqMerge
      -- CP-element group 396: 	 branch_block_stmt_33/forx_xend404x_xloopexit_forx_xend404_PhiReq/$entry
      -- CP-element group 396: 	 branch_block_stmt_33/merge_stmt_1304_PhiAck/dummy
      -- CP-element group 396: 	 branch_block_stmt_33/merge_stmt_1304_PhiAck/$exit
      -- CP-element group 396: 	 branch_block_stmt_33/merge_stmt_1304_PhiAck/$entry
      -- CP-element group 396: 	 branch_block_stmt_33/forx_xbody332_forx_xend404x_xloopexit_PhiReq/$exit
      -- CP-element group 396: 	 branch_block_stmt_33/forx_xbody332_forx_xend404x_xloopexit_PhiReq/$entry
      -- CP-element group 396: 	 branch_block_stmt_33/forx_xbody332_forx_xend404x_xloopexit
      -- 
    if_choice_transition_3029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 396_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1298_branch_ack_1, ack => convTranspose_CP_39_elements(396)); -- 
    -- CP-element group 397:  fork  transition  place  input  output  bypass 
    -- CP-element group 397: predecessors 
    -- CP-element group 397: 	395 
    -- CP-element group 397: successors 
    -- CP-element group 397: 	420 
    -- CP-element group 397: 	421 
    -- CP-element group 397:  members (12) 
      -- CP-element group 397: 	 branch_block_stmt_33/forx_xbody332_forx_xbody332_PhiReq/phi_stmt_1170/phi_stmt_1170_sources/type_cast_1173/$entry
      -- CP-element group 397: 	 branch_block_stmt_33/if_stmt_1298_else_link/$exit
      -- CP-element group 397: 	 branch_block_stmt_33/forx_xbody332_forx_xbody332_PhiReq/phi_stmt_1170/phi_stmt_1170_sources/$entry
      -- CP-element group 397: 	 branch_block_stmt_33/forx_xbody332_forx_xbody332_PhiReq/phi_stmt_1170/phi_stmt_1170_sources/type_cast_1173/SplitProtocol/Sample/$entry
      -- CP-element group 397: 	 branch_block_stmt_33/if_stmt_1298_else_link/else_choice_transition
      -- CP-element group 397: 	 branch_block_stmt_33/forx_xbody332_forx_xbody332_PhiReq/phi_stmt_1170/phi_stmt_1170_sources/type_cast_1173/SplitProtocol/Sample/rr
      -- CP-element group 397: 	 branch_block_stmt_33/forx_xbody332_forx_xbody332_PhiReq/phi_stmt_1170/phi_stmt_1170_sources/type_cast_1173/SplitProtocol/$entry
      -- CP-element group 397: 	 branch_block_stmt_33/forx_xbody332_forx_xbody332_PhiReq/$entry
      -- CP-element group 397: 	 branch_block_stmt_33/forx_xbody332_forx_xbody332
      -- CP-element group 397: 	 branch_block_stmt_33/forx_xbody332_forx_xbody332_PhiReq/phi_stmt_1170/phi_stmt_1170_sources/type_cast_1173/SplitProtocol/Update/cr
      -- CP-element group 397: 	 branch_block_stmt_33/forx_xbody332_forx_xbody332_PhiReq/phi_stmt_1170/$entry
      -- CP-element group 397: 	 branch_block_stmt_33/forx_xbody332_forx_xbody332_PhiReq/phi_stmt_1170/phi_stmt_1170_sources/type_cast_1173/SplitProtocol/Update/$entry
      -- 
    else_choice_transition_3033_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 397_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1298_branch_ack_0, ack => convTranspose_CP_39_elements(397)); -- 
    rr_3308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(397), ack => type_cast_1173_inst_req_0); -- 
    cr_3313_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3313_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(397), ack => type_cast_1173_inst_req_1); -- 
    -- CP-element group 398:  merge  branch  transition  place  output  bypass 
    -- CP-element group 398: predecessors 
    -- CP-element group 398: 	165 
    -- CP-element group 398: 	120 
    -- CP-element group 398: successors 
    -- CP-element group 398: 	121 
    -- CP-element group 398: 	122 
    -- CP-element group 398:  members (17) 
      -- CP-element group 398: 	 branch_block_stmt_33/merge_stmt_402__exit__
      -- CP-element group 398: 	 branch_block_stmt_33/assign_stmt_408__entry__
      -- CP-element group 398: 	 branch_block_stmt_33/assign_stmt_408__exit__
      -- CP-element group 398: 	 branch_block_stmt_33/if_stmt_409__entry__
      -- CP-element group 398: 	 branch_block_stmt_33/merge_stmt_402_PhiReqMerge
      -- CP-element group 398: 	 branch_block_stmt_33/assign_stmt_408/$entry
      -- CP-element group 398: 	 branch_block_stmt_33/assign_stmt_408/$exit
      -- CP-element group 398: 	 branch_block_stmt_33/if_stmt_409_dead_link/$entry
      -- CP-element group 398: 	 branch_block_stmt_33/if_stmt_409_eval_test/$entry
      -- CP-element group 398: 	 branch_block_stmt_33/if_stmt_409_eval_test/$exit
      -- CP-element group 398: 	 branch_block_stmt_33/if_stmt_409_eval_test/branch_req
      -- CP-element group 398: 	 branch_block_stmt_33/R_cmp180413_410_place
      -- CP-element group 398: 	 branch_block_stmt_33/if_stmt_409_if_link/$entry
      -- CP-element group 398: 	 branch_block_stmt_33/if_stmt_409_else_link/$entry
      -- CP-element group 398: 	 branch_block_stmt_33/merge_stmt_402_PhiAck/dummy
      -- CP-element group 398: 	 branch_block_stmt_33/merge_stmt_402_PhiAck/$exit
      -- CP-element group 398: 	 branch_block_stmt_33/merge_stmt_402_PhiAck/$entry
      -- 
    branch_req_925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(398), ack => if_stmt_409_branch_req_0); -- 
    convTranspose_CP_39_elements(398) <= OrReduce(convTranspose_CP_39_elements(165) & convTranspose_CP_39_elements(120));
    -- CP-element group 399:  transition  output  delay-element  bypass 
    -- CP-element group 399: predecessors 
    -- CP-element group 399: 	124 
    -- CP-element group 399: successors 
    -- CP-element group 399: 	403 
    -- CP-element group 399:  members (5) 
      -- CP-element group 399: 	 branch_block_stmt_33/bbx_xnph419_forx_xbody_PhiReq/phi_stmt_453/phi_stmt_453_req
      -- CP-element group 399: 	 branch_block_stmt_33/bbx_xnph419_forx_xbody_PhiReq/phi_stmt_453/phi_stmt_453_sources/type_cast_457_konst_delay_trans
      -- CP-element group 399: 	 branch_block_stmt_33/bbx_xnph419_forx_xbody_PhiReq/phi_stmt_453/phi_stmt_453_sources/$exit
      -- CP-element group 399: 	 branch_block_stmt_33/bbx_xnph419_forx_xbody_PhiReq/phi_stmt_453/$exit
      -- CP-element group 399: 	 branch_block_stmt_33/bbx_xnph419_forx_xbody_PhiReq/$exit
      -- 
    phi_stmt_453_req_3081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_453_req_3081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(399), ack => phi_stmt_453_req_0); -- 
    -- Element group convTranspose_CP_39_elements(399) is a control-delay.
    cp_element_399_delay: control_delay_element  generic map(name => " 399_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(124), ack => convTranspose_CP_39_elements(399), clk => clk, reset =>reset);
    -- CP-element group 400:  transition  input  bypass 
    -- CP-element group 400: predecessors 
    -- CP-element group 400: 	166 
    -- CP-element group 400: successors 
    -- CP-element group 400: 	402 
    -- CP-element group 400:  members (2) 
      -- CP-element group 400: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_453/phi_stmt_453_sources/type_cast_459/SplitProtocol/Sample/ra
      -- CP-element group 400: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_453/phi_stmt_453_sources/type_cast_459/SplitProtocol/Sample/$exit
      -- 
    ra_3101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 400_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_459_inst_ack_0, ack => convTranspose_CP_39_elements(400)); -- 
    -- CP-element group 401:  transition  input  bypass 
    -- CP-element group 401: predecessors 
    -- CP-element group 401: 	166 
    -- CP-element group 401: successors 
    -- CP-element group 401: 	402 
    -- CP-element group 401:  members (2) 
      -- CP-element group 401: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_453/phi_stmt_453_sources/type_cast_459/SplitProtocol/Update/ca
      -- CP-element group 401: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_453/phi_stmt_453_sources/type_cast_459/SplitProtocol/Update/$exit
      -- 
    ca_3106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 401_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_459_inst_ack_1, ack => convTranspose_CP_39_elements(401)); -- 
    -- CP-element group 402:  join  transition  output  bypass 
    -- CP-element group 402: predecessors 
    -- CP-element group 402: 	400 
    -- CP-element group 402: 	401 
    -- CP-element group 402: successors 
    -- CP-element group 402: 	403 
    -- CP-element group 402:  members (6) 
      -- CP-element group 402: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_453/phi_stmt_453_req
      -- CP-element group 402: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_453/phi_stmt_453_sources/type_cast_459/SplitProtocol/$exit
      -- CP-element group 402: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_453/phi_stmt_453_sources/type_cast_459/$exit
      -- CP-element group 402: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_453/phi_stmt_453_sources/$exit
      -- CP-element group 402: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_453/$exit
      -- CP-element group 402: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/$exit
      -- 
    phi_stmt_453_req_3107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_453_req_3107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(402), ack => phi_stmt_453_req_1); -- 
    convTranspose_cp_element_group_402: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_402"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(400) & convTranspose_CP_39_elements(401);
      gj_convTranspose_cp_element_group_402 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(402), clk => clk, reset => reset); --
    end block;
    -- CP-element group 403:  merge  transition  place  bypass 
    -- CP-element group 403: predecessors 
    -- CP-element group 403: 	399 
    -- CP-element group 403: 	402 
    -- CP-element group 403: successors 
    -- CP-element group 403: 	404 
    -- CP-element group 403:  members (2) 
      -- CP-element group 403: 	 branch_block_stmt_33/merge_stmt_452_PhiReqMerge
      -- CP-element group 403: 	 branch_block_stmt_33/merge_stmt_452_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(403) <= OrReduce(convTranspose_CP_39_elements(399) & convTranspose_CP_39_elements(402));
    -- CP-element group 404:  fork  transition  place  input  output  bypass 
    -- CP-element group 404: predecessors 
    -- CP-element group 404: 	403 
    -- CP-element group 404: successors 
    -- CP-element group 404: 	163 
    -- CP-element group 404: 	125 
    -- CP-element group 404: 	126 
    -- CP-element group 404: 	128 
    -- CP-element group 404: 	129 
    -- CP-element group 404: 	132 
    -- CP-element group 404: 	136 
    -- CP-element group 404: 	140 
    -- CP-element group 404: 	144 
    -- CP-element group 404: 	148 
    -- CP-element group 404: 	152 
    -- CP-element group 404: 	156 
    -- CP-element group 404: 	160 
    -- CP-element group 404:  members (56) 
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_Update/$entry
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_558_Update/cr
      -- CP-element group 404: 	 branch_block_stmt_33/merge_stmt_452__exit__
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615__entry__
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_522_update_start_
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_594_update_start_
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_558_Update/$entry
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_558_update_start_
      -- CP-element group 404: 	 branch_block_stmt_33/merge_stmt_452_PhiAck/phi_stmt_453_ack
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_540_Update/cr
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_540_Update/$entry
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_540_update_start_
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_504_Update/cr
      -- CP-element group 404: 	 branch_block_stmt_33/merge_stmt_452_PhiAck/$exit
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_update_start_
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_576_Update/cr
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_504_Update/$entry
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_Update/word_access_complete/word_0/cr
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_576_Update/$entry
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_522_Update/cr
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_Update/word_access_complete/word_0/$entry
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_522_Update/$entry
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_594_Update/cr
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_576_update_start_
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_594_Update/$entry
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_Update/word_access_complete/$entry
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/$entry
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/addr_of_466_update_start_
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_index_resized_1
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_index_scaled_1
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_index_computed_1
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_index_resize_1/$entry
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_index_resize_1/$exit
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_index_resize_1/index_resize_req
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_index_resize_1/index_resize_ack
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_index_scale_1/$entry
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_index_scale_1/$exit
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_index_scale_1/scale_rename_req
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_index_scale_1/scale_rename_ack
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_final_index_sum_regn_update_start
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_final_index_sum_regn_Sample/$entry
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_final_index_sum_regn_Sample/req
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_final_index_sum_regn_Update/$entry
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_final_index_sum_regn_Update/req
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/addr_of_466_complete/$entry
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/addr_of_466_complete/req
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_469_sample_start_
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_469_Sample/$entry
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_469_Sample/rr
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_473_update_start_
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_473_Update/$entry
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_473_Update/cr
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_486_update_start_
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_486_Update/$entry
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_486_Update/cr
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_504_update_start_
      -- 
    phi_stmt_453_ack_3112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 404_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_453_ack_0, ack => convTranspose_CP_39_elements(404)); -- 
    cr_1169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => type_cast_558_inst_req_1); -- 
    cr_1141_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1141_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => type_cast_540_inst_req_1); -- 
    cr_1085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => type_cast_504_inst_req_1); -- 
    cr_1197_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1197_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => type_cast_576_inst_req_1); -- 
    cr_1275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => ptr_deref_602_store_0_req_1); -- 
    cr_1113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => type_cast_522_inst_req_1); -- 
    cr_1225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => type_cast_594_inst_req_1); -- 
    req_981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => array_obj_ref_465_index_offset_req_0); -- 
    req_986_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_986_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => array_obj_ref_465_index_offset_req_1); -- 
    req_1001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => addr_of_466_final_reg_req_1); -- 
    rr_1010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => RPIPE_ConvTranspose_input_pipe_469_inst_req_0); -- 
    cr_1029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => type_cast_473_inst_req_1); -- 
    cr_1057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => type_cast_486_inst_req_1); -- 
    -- CP-element group 405:  transition  output  delay-element  bypass 
    -- CP-element group 405: predecessors 
    -- CP-element group 405: 	168 
    -- CP-element group 405: successors 
    -- CP-element group 405: 	409 
    -- CP-element group 405:  members (5) 
      -- CP-element group 405: 	 branch_block_stmt_33/bbx_xnph415_forx_xbody182_PhiReq/$exit
      -- CP-element group 405: 	 branch_block_stmt_33/bbx_xnph415_forx_xbody182_PhiReq/phi_stmt_660/$exit
      -- CP-element group 405: 	 branch_block_stmt_33/bbx_xnph415_forx_xbody182_PhiReq/phi_stmt_660/phi_stmt_660_sources/$exit
      -- CP-element group 405: 	 branch_block_stmt_33/bbx_xnph415_forx_xbody182_PhiReq/phi_stmt_660/phi_stmt_660_sources/type_cast_666_konst_delay_trans
      -- CP-element group 405: 	 branch_block_stmt_33/bbx_xnph415_forx_xbody182_PhiReq/phi_stmt_660/phi_stmt_660_req
      -- 
    phi_stmt_660_req_3135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_660_req_3135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(405), ack => phi_stmt_660_req_1); -- 
    -- Element group convTranspose_CP_39_elements(405) is a control-delay.
    cp_element_405_delay: control_delay_element  generic map(name => " 405_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(168), ack => convTranspose_CP_39_elements(405), clk => clk, reset =>reset);
    -- CP-element group 406:  transition  input  bypass 
    -- CP-element group 406: predecessors 
    -- CP-element group 406: 	210 
    -- CP-element group 406: successors 
    -- CP-element group 406: 	408 
    -- CP-element group 406:  members (2) 
      -- CP-element group 406: 	 branch_block_stmt_33/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_660/phi_stmt_660_sources/type_cast_663/SplitProtocol/Sample/ra
      -- CP-element group 406: 	 branch_block_stmt_33/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_660/phi_stmt_660_sources/type_cast_663/SplitProtocol/Sample/$exit
      -- 
    ra_3155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 406_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_663_inst_ack_0, ack => convTranspose_CP_39_elements(406)); -- 
    -- CP-element group 407:  transition  input  bypass 
    -- CP-element group 407: predecessors 
    -- CP-element group 407: 	210 
    -- CP-element group 407: successors 
    -- CP-element group 407: 	408 
    -- CP-element group 407:  members (2) 
      -- CP-element group 407: 	 branch_block_stmt_33/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_660/phi_stmt_660_sources/type_cast_663/SplitProtocol/Update/$exit
      -- CP-element group 407: 	 branch_block_stmt_33/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_660/phi_stmt_660_sources/type_cast_663/SplitProtocol/Update/ca
      -- 
    ca_3160_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 407_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_663_inst_ack_1, ack => convTranspose_CP_39_elements(407)); -- 
    -- CP-element group 408:  join  transition  output  bypass 
    -- CP-element group 408: predecessors 
    -- CP-element group 408: 	406 
    -- CP-element group 408: 	407 
    -- CP-element group 408: successors 
    -- CP-element group 408: 	409 
    -- CP-element group 408:  members (6) 
      -- CP-element group 408: 	 branch_block_stmt_33/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_660/phi_stmt_660_sources/type_cast_663/$exit
      -- CP-element group 408: 	 branch_block_stmt_33/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_660/phi_stmt_660_sources/type_cast_663/SplitProtocol/$exit
      -- CP-element group 408: 	 branch_block_stmt_33/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_660/phi_stmt_660_sources/$exit
      -- CP-element group 408: 	 branch_block_stmt_33/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_660/$exit
      -- CP-element group 408: 	 branch_block_stmt_33/forx_xbody182_forx_xbody182_PhiReq/$exit
      -- CP-element group 408: 	 branch_block_stmt_33/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_660/phi_stmt_660_req
      -- 
    phi_stmt_660_req_3161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_660_req_3161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(408), ack => phi_stmt_660_req_0); -- 
    convTranspose_cp_element_group_408: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_408"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(406) & convTranspose_CP_39_elements(407);
      gj_convTranspose_cp_element_group_408 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(408), clk => clk, reset => reset); --
    end block;
    -- CP-element group 409:  merge  transition  place  bypass 
    -- CP-element group 409: predecessors 
    -- CP-element group 409: 	405 
    -- CP-element group 409: 	408 
    -- CP-element group 409: successors 
    -- CP-element group 409: 	410 
    -- CP-element group 409:  members (2) 
      -- CP-element group 409: 	 branch_block_stmt_33/merge_stmt_659_PhiReqMerge
      -- CP-element group 409: 	 branch_block_stmt_33/merge_stmt_659_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(409) <= OrReduce(convTranspose_CP_39_elements(405) & convTranspose_CP_39_elements(408));
    -- CP-element group 410:  fork  transition  place  input  output  bypass 
    -- CP-element group 410: predecessors 
    -- CP-element group 410: 	409 
    -- CP-element group 410: successors 
    -- CP-element group 410: 	188 
    -- CP-element group 410: 	192 
    -- CP-element group 410: 	196 
    -- CP-element group 410: 	200 
    -- CP-element group 410: 	204 
    -- CP-element group 410: 	180 
    -- CP-element group 410: 	184 
    -- CP-element group 410: 	207 
    -- CP-element group 410: 	169 
    -- CP-element group 410: 	170 
    -- CP-element group 410: 	172 
    -- CP-element group 410: 	173 
    -- CP-element group 410: 	176 
    -- CP-element group 410:  members (56) 
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_711_Update/cr
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_711_Update/$entry
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_final_index_sum_regn_update_start
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_711_update_start_
      -- CP-element group 410: 	 branch_block_stmt_33/merge_stmt_659__exit__
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822__entry__
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_693_update_start_
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_676_sample_start_
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/addr_of_673_complete/$entry
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_693_Update/$entry
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_680_update_start_
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_final_index_sum_regn_Update/$entry
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_index_scale_1/scale_rename_ack
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_index_scale_1/scale_rename_req
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_680_Update/cr
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_index_scale_1/$exit
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_index_scale_1/$entry
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_680_Update/$entry
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/addr_of_673_complete/req
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_693_Update/cr
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_final_index_sum_regn_Update/req
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_index_resize_1/index_resize_ack
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_index_resize_1/index_resize_req
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_index_resize_1/$exit
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_index_resize_1/$entry
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_index_computed_1
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_index_scaled_1
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_index_resized_1
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/addr_of_673_update_start_
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/$entry
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_final_index_sum_regn_Sample/req
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_676_Sample/rr
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_final_index_sum_regn_Sample/$entry
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_676_Sample/$entry
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_729_update_start_
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_729_Update/$entry
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_729_Update/cr
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_747_update_start_
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_747_Update/$entry
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_747_Update/cr
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_765_update_start_
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_765_Update/$entry
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_765_Update/cr
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_783_update_start_
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_783_Update/$entry
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_783_Update/cr
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_801_update_start_
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_801_Update/$entry
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_801_Update/cr
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_update_start_
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_Update/$entry
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_Update/word_access_complete/$entry
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_Update/word_access_complete/word_0/$entry
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_Update/word_access_complete/word_0/cr
      -- CP-element group 410: 	 branch_block_stmt_33/merge_stmt_659_PhiAck/phi_stmt_660_ack
      -- CP-element group 410: 	 branch_block_stmt_33/merge_stmt_659_PhiAck/$exit
      -- 
    phi_stmt_660_ack_3166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 410_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_660_ack_0, ack => convTranspose_CP_39_elements(410)); -- 
    cr_1444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(410), ack => type_cast_711_inst_req_1); -- 
    cr_1388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(410), ack => type_cast_680_inst_req_1); -- 
    req_1360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(410), ack => addr_of_673_final_reg_req_1); -- 
    cr_1416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(410), ack => type_cast_693_inst_req_1); -- 
    req_1345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(410), ack => array_obj_ref_672_index_offset_req_1); -- 
    req_1340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(410), ack => array_obj_ref_672_index_offset_req_0); -- 
    rr_1369_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1369_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(410), ack => RPIPE_ConvTranspose_input_pipe_676_inst_req_0); -- 
    cr_1472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(410), ack => type_cast_729_inst_req_1); -- 
    cr_1500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(410), ack => type_cast_747_inst_req_1); -- 
    cr_1528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(410), ack => type_cast_765_inst_req_1); -- 
    cr_1556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(410), ack => type_cast_783_inst_req_1); -- 
    cr_1584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(410), ack => type_cast_801_inst_req_1); -- 
    cr_1634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(410), ack => ptr_deref_809_store_0_req_1); -- 
    -- CP-element group 411:  merge  fork  transition  place  output  bypass 
    -- CP-element group 411: predecessors 
    -- CP-element group 411: 	209 
    -- CP-element group 411: 	122 
    -- CP-element group 411: successors 
    -- CP-element group 411: 	211 
    -- CP-element group 411: 	212 
    -- CP-element group 411: 	213 
    -- CP-element group 411: 	214 
    -- CP-element group 411: 	215 
    -- CP-element group 411: 	216 
    -- CP-element group 411:  members (25) 
      -- CP-element group 411: 	 branch_block_stmt_33/merge_stmt_831__exit__
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859__entry__
      -- CP-element group 411: 	 branch_block_stmt_33/merge_stmt_831_PhiReqMerge
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/$entry
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_834_sample_start_
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_834_update_start_
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_834_Sample/$entry
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_834_Sample/rr
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_834_Update/$entry
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_834_Update/cr
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_838_sample_start_
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_838_update_start_
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_838_Sample/$entry
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_838_Sample/rr
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_838_Update/$entry
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_838_Update/cr
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_842_sample_start_
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_842_update_start_
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_842_Sample/$entry
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_842_Sample/rr
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_842_Update/$entry
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_842_Update/cr
      -- CP-element group 411: 	 branch_block_stmt_33/merge_stmt_831_PhiAck/dummy
      -- CP-element group 411: 	 branch_block_stmt_33/merge_stmt_831_PhiAck/$exit
      -- CP-element group 411: 	 branch_block_stmt_33/merge_stmt_831_PhiAck/$entry
      -- 
    rr_1665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(411), ack => type_cast_834_inst_req_0); -- 
    cr_1670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(411), ack => type_cast_834_inst_req_1); -- 
    rr_1679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(411), ack => type_cast_838_inst_req_0); -- 
    cr_1684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(411), ack => type_cast_838_inst_req_1); -- 
    rr_1693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(411), ack => type_cast_842_inst_req_0); -- 
    cr_1698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(411), ack => type_cast_842_inst_req_1); -- 
    convTranspose_CP_39_elements(411) <= OrReduce(convTranspose_CP_39_elements(209) & convTranspose_CP_39_elements(122));
    -- CP-element group 412:  transition  output  delay-element  bypass 
    -- CP-element group 412: predecessors 
    -- CP-element group 412: 	221 
    -- CP-element group 412: successors 
    -- CP-element group 412: 	416 
    -- CP-element group 412:  members (5) 
      -- CP-element group 412: 	 branch_block_stmt_33/bbx_xnph411_forx_xbody252_PhiReq/phi_stmt_904/phi_stmt_904_req
      -- CP-element group 412: 	 branch_block_stmt_33/bbx_xnph411_forx_xbody252_PhiReq/phi_stmt_904/phi_stmt_904_sources/type_cast_908_konst_delay_trans
      -- CP-element group 412: 	 branch_block_stmt_33/bbx_xnph411_forx_xbody252_PhiReq/phi_stmt_904/phi_stmt_904_sources/$exit
      -- CP-element group 412: 	 branch_block_stmt_33/bbx_xnph411_forx_xbody252_PhiReq/phi_stmt_904/$exit
      -- CP-element group 412: 	 branch_block_stmt_33/bbx_xnph411_forx_xbody252_PhiReq/$exit
      -- 
    phi_stmt_904_req_3212_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_904_req_3212_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(412), ack => phi_stmt_904_req_0); -- 
    -- Element group convTranspose_CP_39_elements(412) is a control-delay.
    cp_element_412_delay: control_delay_element  generic map(name => " 412_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(221), ack => convTranspose_CP_39_elements(412), clk => clk, reset =>reset);
    -- CP-element group 413:  transition  input  bypass 
    -- CP-element group 413: predecessors 
    -- CP-element group 413: 	230 
    -- CP-element group 413: successors 
    -- CP-element group 413: 	415 
    -- CP-element group 413:  members (2) 
      -- CP-element group 413: 	 branch_block_stmt_33/forx_xbody252_forx_xbody252_PhiReq/phi_stmt_904/phi_stmt_904_sources/type_cast_910/SplitProtocol/Sample/ra
      -- CP-element group 413: 	 branch_block_stmt_33/forx_xbody252_forx_xbody252_PhiReq/phi_stmt_904/phi_stmt_904_sources/type_cast_910/SplitProtocol/Sample/$exit
      -- 
    ra_3232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 413_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_910_inst_ack_0, ack => convTranspose_CP_39_elements(413)); -- 
    -- CP-element group 414:  transition  input  bypass 
    -- CP-element group 414: predecessors 
    -- CP-element group 414: 	230 
    -- CP-element group 414: successors 
    -- CP-element group 414: 	415 
    -- CP-element group 414:  members (2) 
      -- CP-element group 414: 	 branch_block_stmt_33/forx_xbody252_forx_xbody252_PhiReq/phi_stmt_904/phi_stmt_904_sources/type_cast_910/SplitProtocol/Update/$exit
      -- CP-element group 414: 	 branch_block_stmt_33/forx_xbody252_forx_xbody252_PhiReq/phi_stmt_904/phi_stmt_904_sources/type_cast_910/SplitProtocol/Update/ca
      -- 
    ca_3237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 414_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_910_inst_ack_1, ack => convTranspose_CP_39_elements(414)); -- 
    -- CP-element group 415:  join  transition  output  bypass 
    -- CP-element group 415: predecessors 
    -- CP-element group 415: 	413 
    -- CP-element group 415: 	414 
    -- CP-element group 415: successors 
    -- CP-element group 415: 	416 
    -- CP-element group 415:  members (6) 
      -- CP-element group 415: 	 branch_block_stmt_33/forx_xbody252_forx_xbody252_PhiReq/phi_stmt_904/phi_stmt_904_sources/$exit
      -- CP-element group 415: 	 branch_block_stmt_33/forx_xbody252_forx_xbody252_PhiReq/phi_stmt_904/phi_stmt_904_sources/type_cast_910/$exit
      -- CP-element group 415: 	 branch_block_stmt_33/forx_xbody252_forx_xbody252_PhiReq/phi_stmt_904/phi_stmt_904_sources/type_cast_910/SplitProtocol/$exit
      -- CP-element group 415: 	 branch_block_stmt_33/forx_xbody252_forx_xbody252_PhiReq/phi_stmt_904/phi_stmt_904_req
      -- CP-element group 415: 	 branch_block_stmt_33/forx_xbody252_forx_xbody252_PhiReq/phi_stmt_904/$exit
      -- CP-element group 415: 	 branch_block_stmt_33/forx_xbody252_forx_xbody252_PhiReq/$exit
      -- 
    phi_stmt_904_req_3238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_904_req_3238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(415), ack => phi_stmt_904_req_1); -- 
    convTranspose_cp_element_group_415: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_415"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(413) & convTranspose_CP_39_elements(414);
      gj_convTranspose_cp_element_group_415 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(415), clk => clk, reset => reset); --
    end block;
    -- CP-element group 416:  merge  transition  place  bypass 
    -- CP-element group 416: predecessors 
    -- CP-element group 416: 	412 
    -- CP-element group 416: 	415 
    -- CP-element group 416: successors 
    -- CP-element group 416: 	417 
    -- CP-element group 416:  members (2) 
      -- CP-element group 416: 	 branch_block_stmt_33/merge_stmt_903_PhiReqMerge
      -- CP-element group 416: 	 branch_block_stmt_33/merge_stmt_903_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(416) <= OrReduce(convTranspose_CP_39_elements(412) & convTranspose_CP_39_elements(415));
    -- CP-element group 417:  fork  transition  place  input  output  bypass 
    -- CP-element group 417: predecessors 
    -- CP-element group 417: 	416 
    -- CP-element group 417: successors 
    -- CP-element group 417: 	222 
    -- CP-element group 417: 	223 
    -- CP-element group 417: 	225 
    -- CP-element group 417: 	227 
    -- CP-element group 417:  members (29) 
      -- CP-element group 417: 	 branch_block_stmt_33/merge_stmt_903__exit__
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934__entry__
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/$entry
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/addr_of_917_update_start_
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_index_resized_1
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_index_scaled_1
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_index_computed_1
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_index_resize_1/$entry
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_index_resize_1/$exit
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_index_resize_1/index_resize_req
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_index_resize_1/index_resize_ack
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_index_scale_1/$entry
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_index_scale_1/$exit
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_index_scale_1/scale_rename_req
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_index_scale_1/scale_rename_ack
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_final_index_sum_regn_update_start
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_final_index_sum_regn_Sample/$entry
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_final_index_sum_regn_Sample/req
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_final_index_sum_regn_Update/$entry
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_final_index_sum_regn_Update/req
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/addr_of_917_complete/$entry
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/addr_of_917_complete/req
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_update_start_
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_Update/$entry
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_Update/word_access_complete/$entry
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_Update/word_access_complete/word_0/$entry
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_Update/word_access_complete/word_0/cr
      -- CP-element group 417: 	 branch_block_stmt_33/merge_stmt_903_PhiAck/phi_stmt_904_ack
      -- CP-element group 417: 	 branch_block_stmt_33/merge_stmt_903_PhiAck/$exit
      -- 
    phi_stmt_904_ack_3243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 417_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_904_ack_0, ack => convTranspose_CP_39_elements(417)); -- 
    req_1763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(417), ack => array_obj_ref_916_index_offset_req_0); -- 
    req_1768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(417), ack => array_obj_ref_916_index_offset_req_1); -- 
    req_1783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(417), ack => addr_of_917_final_reg_req_1); -- 
    cr_1833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(417), ack => ptr_deref_920_store_0_req_1); -- 
    -- CP-element group 418:  merge  fork  transition  place  output  bypass 
    -- CP-element group 418: predecessors 
    -- CP-element group 418: 	219 
    -- CP-element group 418: 	229 
    -- CP-element group 418: successors 
    -- CP-element group 418: 	283 
    -- CP-element group 418: 	307 
    -- CP-element group 418: 	331 
    -- CP-element group 418: 	333 
    -- CP-element group 418: 	335 
    -- CP-element group 418: 	337 
    -- CP-element group 418: 	231 
    -- CP-element group 418: 	232 
    -- CP-element group 418: 	234 
    -- CP-element group 418: 	235 
    -- CP-element group 418: 	259 
    -- CP-element group 418:  members (40) 
      -- CP-element group 418: 	 branch_block_stmt_33/merge_stmt_943__exit__
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108__entry__
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1061_Sample/req
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1061_Sample/$entry
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1061_sample_start_
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1025_Sample/req
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1025_Sample/$entry
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_989_Sample/req
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_989_Sample/$entry
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_989_sample_start_
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1025_sample_start_
      -- CP-element group 418: 	 branch_block_stmt_33/merge_stmt_943_PhiReqMerge
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/$entry
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/call_stmt_946_sample_start_
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/call_stmt_946_update_start_
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/call_stmt_946_Sample/$entry
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/call_stmt_946_Sample/crr
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/call_stmt_946_Update/$entry
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/call_stmt_946_Update/ccr
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/type_cast_951_update_start_
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/type_cast_951_Update/$entry
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/type_cast_951_Update/cr
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_953_sample_start_
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_953_Sample/$entry
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_953_Sample/req
      -- CP-element group 418: 	 branch_block_stmt_33/merge_stmt_943_PhiAck/dummy
      -- CP-element group 418: 	 branch_block_stmt_33/merge_stmt_943_PhiAck/$exit
      -- CP-element group 418: 	 branch_block_stmt_33/merge_stmt_943_PhiAck/$entry
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block0_done_1098_sample_start_
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block0_done_1098_Sample/$entry
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block0_done_1098_Sample/rr
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block1_done_1101_sample_start_
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block1_done_1101_Sample/$entry
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block1_done_1101_Sample/rr
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block2_done_1104_sample_start_
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block2_done_1104_Sample/$entry
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block2_done_1104_Sample/rr
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block3_done_1107_sample_start_
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block3_done_1107_Sample/$entry
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block3_done_1107_Sample/rr
      -- 
    req_2396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(418), ack => WPIPE_Block3_start_1061_inst_req_0); -- 
    req_2228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(418), ack => WPIPE_Block2_start_1025_inst_req_0); -- 
    req_2060_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2060_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(418), ack => WPIPE_Block1_start_989_inst_req_0); -- 
    crr_1864_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1864_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(418), ack => call_stmt_946_call_req_0); -- 
    ccr_1869_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1869_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(418), ack => call_stmt_946_call_req_1); -- 
    cr_1883_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1883_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(418), ack => type_cast_951_inst_req_1); -- 
    req_1892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(418), ack => WPIPE_Block0_start_953_inst_req_0); -- 
    rr_2564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(418), ack => RPIPE_Block0_done_1098_inst_req_0); -- 
    rr_2578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(418), ack => RPIPE_Block1_done_1101_inst_req_0); -- 
    rr_2592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(418), ack => RPIPE_Block2_done_1104_inst_req_0); -- 
    rr_2606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(418), ack => RPIPE_Block3_done_1107_inst_req_0); -- 
    convTranspose_CP_39_elements(418) <= OrReduce(convTranspose_CP_39_elements(219) & convTranspose_CP_39_elements(229));
    -- CP-element group 419:  transition  output  delay-element  bypass 
    -- CP-element group 419: predecessors 
    -- CP-element group 419: 	349 
    -- CP-element group 419: successors 
    -- CP-element group 419: 	423 
    -- CP-element group 419:  members (5) 
      -- CP-element group 419: 	 branch_block_stmt_33/bbx_xnph_forx_xbody332_PhiReq/$exit
      -- CP-element group 419: 	 branch_block_stmt_33/bbx_xnph_forx_xbody332_PhiReq/phi_stmt_1170/$exit
      -- CP-element group 419: 	 branch_block_stmt_33/bbx_xnph_forx_xbody332_PhiReq/phi_stmt_1170/phi_stmt_1170_sources/$exit
      -- CP-element group 419: 	 branch_block_stmt_33/bbx_xnph_forx_xbody332_PhiReq/phi_stmt_1170/phi_stmt_1170_sources/type_cast_1176_konst_delay_trans
      -- CP-element group 419: 	 branch_block_stmt_33/bbx_xnph_forx_xbody332_PhiReq/phi_stmt_1170/phi_stmt_1170_req
      -- 
    phi_stmt_1170_req_3289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1170_req_3289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(419), ack => phi_stmt_1170_req_1); -- 
    -- Element group convTranspose_CP_39_elements(419) is a control-delay.
    cp_element_419_delay: control_delay_element  generic map(name => " 419_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(349), ack => convTranspose_CP_39_elements(419), clk => clk, reset =>reset);
    -- CP-element group 420:  transition  input  bypass 
    -- CP-element group 420: predecessors 
    -- CP-element group 420: 	397 
    -- CP-element group 420: successors 
    -- CP-element group 420: 	422 
    -- CP-element group 420:  members (2) 
      -- CP-element group 420: 	 branch_block_stmt_33/forx_xbody332_forx_xbody332_PhiReq/phi_stmt_1170/phi_stmt_1170_sources/type_cast_1173/SplitProtocol/Sample/$exit
      -- CP-element group 420: 	 branch_block_stmt_33/forx_xbody332_forx_xbody332_PhiReq/phi_stmt_1170/phi_stmt_1170_sources/type_cast_1173/SplitProtocol/Sample/ra
      -- 
    ra_3309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 420_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1173_inst_ack_0, ack => convTranspose_CP_39_elements(420)); -- 
    -- CP-element group 421:  transition  input  bypass 
    -- CP-element group 421: predecessors 
    -- CP-element group 421: 	397 
    -- CP-element group 421: successors 
    -- CP-element group 421: 	422 
    -- CP-element group 421:  members (2) 
      -- CP-element group 421: 	 branch_block_stmt_33/forx_xbody332_forx_xbody332_PhiReq/phi_stmt_1170/phi_stmt_1170_sources/type_cast_1173/SplitProtocol/Update/ca
      -- CP-element group 421: 	 branch_block_stmt_33/forx_xbody332_forx_xbody332_PhiReq/phi_stmt_1170/phi_stmt_1170_sources/type_cast_1173/SplitProtocol/Update/$exit
      -- 
    ca_3314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 421_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1173_inst_ack_1, ack => convTranspose_CP_39_elements(421)); -- 
    -- CP-element group 422:  join  transition  output  bypass 
    -- CP-element group 422: predecessors 
    -- CP-element group 422: 	420 
    -- CP-element group 422: 	421 
    -- CP-element group 422: successors 
    -- CP-element group 422: 	423 
    -- CP-element group 422:  members (6) 
      -- CP-element group 422: 	 branch_block_stmt_33/forx_xbody332_forx_xbody332_PhiReq/$exit
      -- CP-element group 422: 	 branch_block_stmt_33/forx_xbody332_forx_xbody332_PhiReq/phi_stmt_1170/phi_stmt_1170_sources/type_cast_1173/SplitProtocol/$exit
      -- CP-element group 422: 	 branch_block_stmt_33/forx_xbody332_forx_xbody332_PhiReq/phi_stmt_1170/phi_stmt_1170_sources/$exit
      -- CP-element group 422: 	 branch_block_stmt_33/forx_xbody332_forx_xbody332_PhiReq/phi_stmt_1170/phi_stmt_1170_sources/type_cast_1173/$exit
      -- CP-element group 422: 	 branch_block_stmt_33/forx_xbody332_forx_xbody332_PhiReq/phi_stmt_1170/phi_stmt_1170_req
      -- CP-element group 422: 	 branch_block_stmt_33/forx_xbody332_forx_xbody332_PhiReq/phi_stmt_1170/$exit
      -- 
    phi_stmt_1170_req_3315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1170_req_3315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(422), ack => phi_stmt_1170_req_0); -- 
    convTranspose_cp_element_group_422: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_422"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(420) & convTranspose_CP_39_elements(421);
      gj_convTranspose_cp_element_group_422 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(422), clk => clk, reset => reset); --
    end block;
    -- CP-element group 423:  merge  transition  place  bypass 
    -- CP-element group 423: predecessors 
    -- CP-element group 423: 	419 
    -- CP-element group 423: 	422 
    -- CP-element group 423: successors 
    -- CP-element group 423: 	424 
    -- CP-element group 423:  members (2) 
      -- CP-element group 423: 	 branch_block_stmt_33/merge_stmt_1169_PhiReqMerge
      -- CP-element group 423: 	 branch_block_stmt_33/merge_stmt_1169_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(423) <= OrReduce(convTranspose_CP_39_elements(419) & convTranspose_CP_39_elements(422));
    -- CP-element group 424:  fork  transition  place  input  output  bypass 
    -- CP-element group 424: predecessors 
    -- CP-element group 424: 	423 
    -- CP-element group 424: successors 
    -- CP-element group 424: 	350 
    -- CP-element group 424: 	351 
    -- CP-element group 424: 	353 
    -- CP-element group 424: 	355 
    -- CP-element group 424: 	357 
    -- CP-element group 424: 	359 
    -- CP-element group 424: 	361 
    -- CP-element group 424: 	363 
    -- CP-element group 424: 	365 
    -- CP-element group 424: 	367 
    -- CP-element group 424: 	369 
    -- CP-element group 424: 	371 
    -- CP-element group 424:  members (53) 
      -- CP-element group 424: 	 branch_block_stmt_33/merge_stmt_1169__exit__
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297__entry__
      -- CP-element group 424: 	 branch_block_stmt_33/merge_stmt_1169_PhiAck/$exit
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/$entry
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/addr_of_1183_update_start_
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/array_obj_ref_1182_index_resized_1
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/array_obj_ref_1182_index_scaled_1
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/array_obj_ref_1182_index_computed_1
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/array_obj_ref_1182_index_resize_1/$entry
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/array_obj_ref_1182_index_resize_1/$exit
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/array_obj_ref_1182_index_resize_1/index_resize_req
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/array_obj_ref_1182_index_resize_1/index_resize_ack
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/array_obj_ref_1182_index_scale_1/$entry
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/array_obj_ref_1182_index_scale_1/$exit
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/array_obj_ref_1182_index_scale_1/scale_rename_req
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/array_obj_ref_1182_index_scale_1/scale_rename_ack
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/array_obj_ref_1182_final_index_sum_regn_update_start
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/array_obj_ref_1182_final_index_sum_regn_Sample/$entry
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/array_obj_ref_1182_final_index_sum_regn_Sample/req
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/array_obj_ref_1182_final_index_sum_regn_Update/$entry
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/array_obj_ref_1182_final_index_sum_regn_Update/req
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/addr_of_1183_complete/$entry
      -- CP-element group 424: 	 branch_block_stmt_33/merge_stmt_1169_PhiAck/phi_stmt_1170_ack
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/addr_of_1183_complete/req
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/ptr_deref_1187_update_start_
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/ptr_deref_1187_Update/$entry
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/ptr_deref_1187_Update/word_access_complete/$entry
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/ptr_deref_1187_Update/word_access_complete/word_0/$entry
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/ptr_deref_1187_Update/word_access_complete/word_0/cr
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1191_update_start_
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1191_Update/$entry
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1191_Update/cr
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1201_update_start_
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1201_Update/$entry
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1201_Update/cr
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1211_update_start_
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1211_Update/$entry
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1211_Update/cr
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1221_update_start_
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1221_Update/$entry
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1221_Update/cr
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1231_update_start_
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1231_Update/$entry
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1231_Update/cr
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1241_update_start_
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1241_Update/$entry
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1241_Update/cr
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1251_update_start_
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1251_Update/$entry
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1251_Update/cr
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1261_update_start_
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1261_Update/$entry
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1184_to_assign_stmt_1297/type_cast_1261_Update/cr
      -- 
    phi_stmt_1170_ack_3320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 424_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1170_ack_0, ack => convTranspose_CP_39_elements(424)); -- 
    req_2721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(424), ack => array_obj_ref_1182_index_offset_req_0); -- 
    req_2726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(424), ack => array_obj_ref_1182_index_offset_req_1); -- 
    req_2741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(424), ack => addr_of_1183_final_reg_req_1); -- 
    cr_2786_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2786_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(424), ack => ptr_deref_1187_load_0_req_1); -- 
    cr_2805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(424), ack => type_cast_1191_inst_req_1); -- 
    cr_2819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(424), ack => type_cast_1201_inst_req_1); -- 
    cr_2833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(424), ack => type_cast_1211_inst_req_1); -- 
    cr_2847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(424), ack => type_cast_1221_inst_req_1); -- 
    cr_2861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(424), ack => type_cast_1231_inst_req_1); -- 
    cr_2875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(424), ack => type_cast_1241_inst_req_1); -- 
    cr_2889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(424), ack => type_cast_1251_inst_req_1); -- 
    cr_2903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(424), ack => type_cast_1261_inst_req_1); -- 
    -- CP-element group 425:  merge  transition  place  bypass 
    -- CP-element group 425: predecessors 
    -- CP-element group 425: 	347 
    -- CP-element group 425: 	396 
    -- CP-element group 425: successors 
    -- CP-element group 425:  members (16) 
      -- CP-element group 425: 	 $exit
      -- CP-element group 425: 	 branch_block_stmt_33/$exit
      -- CP-element group 425: 	 branch_block_stmt_33/branch_block_stmt_33__exit__
      -- CP-element group 425: 	 branch_block_stmt_33/merge_stmt_1306__exit__
      -- CP-element group 425: 	 branch_block_stmt_33/return__
      -- CP-element group 425: 	 branch_block_stmt_33/merge_stmt_1308__exit__
      -- CP-element group 425: 	 branch_block_stmt_33/merge_stmt_1306_PhiAck/$exit
      -- CP-element group 425: 	 branch_block_stmt_33/merge_stmt_1306_PhiAck/$entry
      -- CP-element group 425: 	 branch_block_stmt_33/merge_stmt_1306_PhiAck/dummy
      -- CP-element group 425: 	 branch_block_stmt_33/return___PhiReq/$entry
      -- CP-element group 425: 	 branch_block_stmt_33/return___PhiReq/$exit
      -- CP-element group 425: 	 branch_block_stmt_33/merge_stmt_1306_PhiReqMerge
      -- CP-element group 425: 	 branch_block_stmt_33/merge_stmt_1308_PhiReqMerge
      -- CP-element group 425: 	 branch_block_stmt_33/merge_stmt_1308_PhiAck/$entry
      -- CP-element group 425: 	 branch_block_stmt_33/merge_stmt_1308_PhiAck/dummy
      -- CP-element group 425: 	 branch_block_stmt_33/merge_stmt_1308_PhiAck/$exit
      -- 
    convTranspose_CP_39_elements(425) <= OrReduce(convTranspose_CP_39_elements(347) & convTranspose_CP_39_elements(396));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar429_915_resized : std_logic_vector(13 downto 0);
    signal R_indvar429_915_scaled : std_logic_vector(13 downto 0);
    signal R_indvar443_671_resized : std_logic_vector(10 downto 0);
    signal R_indvar443_671_scaled : std_logic_vector(10 downto 0);
    signal R_indvar459_464_resized : std_logic_vector(13 downto 0);
    signal R_indvar459_464_scaled : std_logic_vector(13 downto 0);
    signal R_indvar_1181_resized : std_logic_vector(13 downto 0);
    signal R_indvar_1181_scaled : std_logic_vector(13 downto 0);
    signal add104_336 : std_logic_vector(15 downto 0);
    signal add113_361 : std_logic_vector(15 downto 0);
    signal add122_386 : std_logic_vector(15 downto 0);
    signal add12_83 : std_logic_vector(15 downto 0);
    signal add136_492 : std_logic_vector(63 downto 0);
    signal add142_510 : std_logic_vector(63 downto 0);
    signal add148_528 : std_logic_vector(63 downto 0);
    signal add154_546 : std_logic_vector(63 downto 0);
    signal add160_564 : std_logic_vector(63 downto 0);
    signal add166_582 : std_logic_vector(63 downto 0);
    signal add172_600 : std_logic_vector(63 downto 0);
    signal add192_699 : std_logic_vector(63 downto 0);
    signal add198_717 : std_logic_vector(63 downto 0);
    signal add204_735 : std_logic_vector(63 downto 0);
    signal add210_753 : std_logic_vector(63 downto 0);
    signal add216_771 : std_logic_vector(63 downto 0);
    signal add21_108 : std_logic_vector(15 downto 0);
    signal add222_789 : std_logic_vector(63 downto 0);
    signal add228_807 : std_logic_vector(63 downto 0);
    signal add30_133 : std_logic_vector(15 downto 0);
    signal add39_158 : std_logic_vector(15 downto 0);
    signal add48_183 : std_logic_vector(15 downto 0);
    signal add57_208 : std_logic_vector(15 downto 0);
    signal add86_286 : std_logic_vector(15 downto 0);
    signal add95_311 : std_logic_vector(15 downto 0);
    signal add_58 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1182_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1182_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1182_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1182_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1182_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1182_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_465_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_465_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_465_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_465_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_465_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_465_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_672_constant_part_of_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_672_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_672_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_672_offset_scale_factor_1 : std_logic_vector(10 downto 0);
    signal array_obj_ref_672_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_672_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_916_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_916_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_916_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_916_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_916_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_916_root_address : std_logic_vector(13 downto 0);
    signal arrayidx232_674 : std_logic_vector(31 downto 0);
    signal arrayidx255_918 : std_logic_vector(31 downto 0);
    signal arrayidx337_1184 : std_logic_vector(31 downto 0);
    signal arrayidx_467 : std_logic_vector(31 downto 0);
    signal call102_327 : std_logic_vector(7 downto 0);
    signal call106_339 : std_logic_vector(7 downto 0);
    signal call10_74 : std_logic_vector(7 downto 0);
    signal call111_352 : std_logic_vector(7 downto 0);
    signal call115_364 : std_logic_vector(7 downto 0);
    signal call120_377 : std_logic_vector(7 downto 0);
    signal call129_470 : std_logic_vector(7 downto 0);
    signal call133_483 : std_logic_vector(7 downto 0);
    signal call139_501 : std_logic_vector(7 downto 0);
    signal call145_519 : std_logic_vector(7 downto 0);
    signal call14_86 : std_logic_vector(7 downto 0);
    signal call151_537 : std_logic_vector(7 downto 0);
    signal call157_555 : std_logic_vector(7 downto 0);
    signal call163_573 : std_logic_vector(7 downto 0);
    signal call169_591 : std_logic_vector(7 downto 0);
    signal call185_677 : std_logic_vector(7 downto 0);
    signal call189_690 : std_logic_vector(7 downto 0);
    signal call195_708 : std_logic_vector(7 downto 0);
    signal call19_99 : std_logic_vector(7 downto 0);
    signal call201_726 : std_logic_vector(7 downto 0);
    signal call207_744 : std_logic_vector(7 downto 0);
    signal call213_762 : std_logic_vector(7 downto 0);
    signal call219_780 : std_logic_vector(7 downto 0);
    signal call225_798 : std_logic_vector(7 downto 0);
    signal call23_111 : std_logic_vector(7 downto 0);
    signal call261_946 : std_logic_vector(63 downto 0);
    signal call28_124 : std_logic_vector(7 downto 0);
    signal call2_49 : std_logic_vector(7 downto 0);
    signal call312_1099 : std_logic_vector(15 downto 0);
    signal call314_1102 : std_logic_vector(15 downto 0);
    signal call316_1105 : std_logic_vector(15 downto 0);
    signal call318_1108 : std_logic_vector(15 downto 0);
    signal call320_1111 : std_logic_vector(63 downto 0);
    signal call32_136 : std_logic_vector(7 downto 0);
    signal call37_149 : std_logic_vector(7 downto 0);
    signal call41_161 : std_logic_vector(7 downto 0);
    signal call46_174 : std_logic_vector(7 downto 0);
    signal call50_186 : std_logic_vector(7 downto 0);
    signal call55_199 : std_logic_vector(7 downto 0);
    signal call5_61 : std_logic_vector(7 downto 0);
    signal call79_264 : std_logic_vector(7 downto 0);
    signal call84_277 : std_logic_vector(7 downto 0);
    signal call88_289 : std_logic_vector(7 downto 0);
    signal call93_302 : std_logic_vector(7 downto 0);
    signal call97_314 : std_logic_vector(7 downto 0);
    signal call_36 : std_logic_vector(7 downto 0);
    signal cmp180413_408 : std_logic_vector(0 downto 0);
    signal cmp250409_859 : std_logic_vector(0 downto 0);
    signal cmp417_393 : std_logic_vector(0 downto 0);
    signal conv100_318 : std_logic_vector(15 downto 0);
    signal conv103_331 : std_logic_vector(15 downto 0);
    signal conv109_343 : std_logic_vector(15 downto 0);
    signal conv112_356 : std_logic_vector(15 downto 0);
    signal conv118_368 : std_logic_vector(15 downto 0);
    signal conv11_78 : std_logic_vector(15 downto 0);
    signal conv121_381 : std_logic_vector(15 downto 0);
    signal conv130_474 : std_logic_vector(63 downto 0);
    signal conv135_487 : std_logic_vector(63 downto 0);
    signal conv141_505 : std_logic_vector(63 downto 0);
    signal conv147_523 : std_logic_vector(63 downto 0);
    signal conv153_541 : std_logic_vector(63 downto 0);
    signal conv159_559 : std_logic_vector(63 downto 0);
    signal conv165_577 : std_logic_vector(63 downto 0);
    signal conv171_595 : std_logic_vector(63 downto 0);
    signal conv17_90 : std_logic_vector(15 downto 0);
    signal conv186_681 : std_logic_vector(63 downto 0);
    signal conv191_694 : std_logic_vector(63 downto 0);
    signal conv197_712 : std_logic_vector(63 downto 0);
    signal conv1_40 : std_logic_vector(15 downto 0);
    signal conv203_730 : std_logic_vector(63 downto 0);
    signal conv209_748 : std_logic_vector(63 downto 0);
    signal conv20_103 : std_logic_vector(15 downto 0);
    signal conv215_766 : std_logic_vector(63 downto 0);
    signal conv221_784 : std_logic_vector(63 downto 0);
    signal conv227_802 : std_logic_vector(63 downto 0);
    signal conv239_835 : std_logic_vector(31 downto 0);
    signal conv241_839 : std_logic_vector(31 downto 0);
    signal conv244_843 : std_logic_vector(31 downto 0);
    signal conv262_952 : std_logic_vector(63 downto 0);
    signal conv26_115 : std_logic_vector(15 downto 0);
    signal conv29_128 : std_logic_vector(15 downto 0);
    signal conv321_1116 : std_logic_vector(63 downto 0);
    signal conv341_1192 : std_logic_vector(7 downto 0);
    signal conv347_1202 : std_logic_vector(7 downto 0);
    signal conv353_1212 : std_logic_vector(7 downto 0);
    signal conv359_1222 : std_logic_vector(7 downto 0);
    signal conv35_140 : std_logic_vector(15 downto 0);
    signal conv365_1232 : std_logic_vector(7 downto 0);
    signal conv371_1242 : std_logic_vector(7 downto 0);
    signal conv377_1252 : std_logic_vector(7 downto 0);
    signal conv383_1262 : std_logic_vector(7 downto 0);
    signal conv38_153 : std_logic_vector(15 downto 0);
    signal conv3_53 : std_logic_vector(15 downto 0);
    signal conv44_165 : std_logic_vector(15 downto 0);
    signal conv47_178 : std_logic_vector(15 downto 0);
    signal conv53_190 : std_logic_vector(15 downto 0);
    signal conv56_203 : std_logic_vector(15 downto 0);
    signal conv61_212 : std_logic_vector(31 downto 0);
    signal conv63_216 : std_logic_vector(31 downto 0);
    signal conv65_220 : std_logic_vector(31 downto 0);
    signal conv69_234 : std_logic_vector(31 downto 0);
    signal conv71_238 : std_logic_vector(31 downto 0);
    signal conv74_242 : std_logic_vector(31 downto 0);
    signal conv77_246 : std_logic_vector(31 downto 0);
    signal conv82_268 : std_logic_vector(15 downto 0);
    signal conv85_281 : std_logic_vector(15 downto 0);
    signal conv8_65 : std_logic_vector(15 downto 0);
    signal conv91_293 : std_logic_vector(15 downto 0);
    signal conv94_306 : std_logic_vector(15 downto 0);
    signal exitcond1_1297 : std_logic_vector(0 downto 0);
    signal exitcond2_822 : std_logic_vector(0 downto 0);
    signal exitcond3_615 : std_logic_vector(0 downto 0);
    signal exitcond_934 : std_logic_vector(0 downto 0);
    signal iNsTr_163_1154 : std_logic_vector(63 downto 0);
    signal iNsTr_25_437 : std_logic_vector(63 downto 0);
    signal iNsTr_38_644 : std_logic_vector(63 downto 0);
    signal iNsTr_52_888 : std_logic_vector(63 downto 0);
    signal indvar429_904 : std_logic_vector(63 downto 0);
    signal indvar443_660 : std_logic_vector(63 downto 0);
    signal indvar459_453 : std_logic_vector(63 downto 0);
    signal indvar_1170 : std_logic_vector(63 downto 0);
    signal indvarx_xnext430_929 : std_logic_vector(63 downto 0);
    signal indvarx_xnext444_817 : std_logic_vector(63 downto 0);
    signal indvarx_xnext460_610 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1292 : std_logic_vector(63 downto 0);
    signal mul242_848 : std_logic_vector(31 downto 0);
    signal mul245_853 : std_logic_vector(31 downto 0);
    signal mul66_230 : std_logic_vector(31 downto 0);
    signal mul72_251 : std_logic_vector(31 downto 0);
    signal mul75_256 : std_logic_vector(31 downto 0);
    signal mul78_261 : std_logic_vector(31 downto 0);
    signal mul_225 : std_logic_vector(31 downto 0);
    signal ptr_deref_1187_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1187_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1187_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1187_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1187_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_602_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_602_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_602_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_602_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_602_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_602_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_809_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_809_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_809_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_809_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_809_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_809_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_920_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_920_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_920_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_920_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_920_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_920_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl101_324 : std_logic_vector(15 downto 0);
    signal shl110_349 : std_logic_vector(15 downto 0);
    signal shl119_374 : std_logic_vector(15 downto 0);
    signal shl132_480 : std_logic_vector(63 downto 0);
    signal shl138_498 : std_logic_vector(63 downto 0);
    signal shl144_516 : std_logic_vector(63 downto 0);
    signal shl150_534 : std_logic_vector(63 downto 0);
    signal shl156_552 : std_logic_vector(63 downto 0);
    signal shl162_570 : std_logic_vector(63 downto 0);
    signal shl168_588 : std_logic_vector(63 downto 0);
    signal shl188_687 : std_logic_vector(63 downto 0);
    signal shl18_96 : std_logic_vector(15 downto 0);
    signal shl194_705 : std_logic_vector(63 downto 0);
    signal shl200_723 : std_logic_vector(63 downto 0);
    signal shl206_741 : std_logic_vector(63 downto 0);
    signal shl212_759 : std_logic_vector(63 downto 0);
    signal shl218_777 : std_logic_vector(63 downto 0);
    signal shl224_795 : std_logic_vector(63 downto 0);
    signal shl27_121 : std_logic_vector(15 downto 0);
    signal shl36_146 : std_logic_vector(15 downto 0);
    signal shl45_171 : std_logic_vector(15 downto 0);
    signal shl54_196 : std_logic_vector(15 downto 0);
    signal shl83_274 : std_logic_vector(15 downto 0);
    signal shl92_299 : std_logic_vector(15 downto 0);
    signal shl9_71 : std_logic_vector(15 downto 0);
    signal shl_46 : std_logic_vector(15 downto 0);
    signal shr344_1198 : std_logic_vector(63 downto 0);
    signal shr350_1208 : std_logic_vector(63 downto 0);
    signal shr356_1218 : std_logic_vector(63 downto 0);
    signal shr362_1228 : std_logic_vector(63 downto 0);
    signal shr368_1238 : std_logic_vector(63 downto 0);
    signal shr374_1248 : std_logic_vector(63 downto 0);
    signal shr380_1258 : std_logic_vector(63 downto 0);
    signal sub_1121 : std_logic_vector(63 downto 0);
    signal tmp338_1188 : std_logic_vector(63 downto 0);
    signal tmp424_1138 : std_logic_vector(31 downto 0);
    signal tmp424x_xop_1150 : std_logic_vector(31 downto 0);
    signal tmp425_1144 : std_logic_vector(0 downto 0);
    signal tmp428_1167 : std_logic_vector(63 downto 0);
    signal tmp436_872 : std_logic_vector(31 downto 0);
    signal tmp436x_xop_884 : std_logic_vector(31 downto 0);
    signal tmp437_878 : std_logic_vector(0 downto 0);
    signal tmp441_901 : std_logic_vector(63 downto 0);
    signal tmp452_628 : std_logic_vector(31 downto 0);
    signal tmp452x_xop_640 : std_logic_vector(31 downto 0);
    signal tmp453_634 : std_logic_vector(0 downto 0);
    signal tmp457_657 : std_logic_vector(63 downto 0);
    signal tmp466_421 : std_logic_vector(31 downto 0);
    signal tmp466x_xop_433 : std_logic_vector(31 downto 0);
    signal tmp467_427 : std_logic_vector(0 downto 0);
    signal tmp471_450 : std_logic_vector(63 downto 0);
    signal type_cast_1114_wire : std_logic_vector(63 downto 0);
    signal type_cast_1136_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1142_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1148_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1158_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1165_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1173_wire : std_logic_vector(63 downto 0);
    signal type_cast_1176_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1196_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_119_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1206_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1216_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1226_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1236_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1246_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1256_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1290_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_144_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_169_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_194_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_272_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_297_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_322_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_347_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_372_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_390_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_406_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_419_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_425_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_431_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_441_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_448_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_44_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_457_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_459_wire : std_logic_vector(63 downto 0);
    signal type_cast_478_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_496_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_514_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_532_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_550_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_568_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_586_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_608_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_626_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_632_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_638_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_648_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_655_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_663_wire : std_logic_vector(63 downto 0);
    signal type_cast_666_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_685_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_69_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_703_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_721_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_739_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_757_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_775_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_793_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_815_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_857_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_870_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_876_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_882_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_892_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_899_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_908_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_910_wire : std_logic_vector(63 downto 0);
    signal type_cast_922_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_927_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_94_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_950_wire : std_logic_vector(63 downto 0);
    signal xx_xop473_894 : std_logic_vector(63 downto 0);
    signal xx_xop474_650 : std_logic_vector(63 downto 0);
    signal xx_xop475_443 : std_logic_vector(63 downto 0);
    signal xx_xop_1160 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1182_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1182_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1182_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1182_resized_base_address <= "00000000000000";
    array_obj_ref_465_constant_part_of_offset <= "00000000000000";
    array_obj_ref_465_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_465_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_465_resized_base_address <= "00000000000000";
    array_obj_ref_672_constant_part_of_offset <= "00000100010";
    array_obj_ref_672_offset_scale_factor_0 <= "10000000000";
    array_obj_ref_672_offset_scale_factor_1 <= "00000000001";
    array_obj_ref_672_resized_base_address <= "00000000000";
    array_obj_ref_916_constant_part_of_offset <= "00000000000000";
    array_obj_ref_916_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_916_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_916_resized_base_address <= "00000000000000";
    ptr_deref_1187_word_offset_0 <= "00000000000000";
    ptr_deref_602_word_offset_0 <= "00000000000000";
    ptr_deref_809_word_offset_0 <= "00000000000";
    ptr_deref_920_word_offset_0 <= "00000000000000";
    type_cast_1136_wire_constant <= "00000000000000000000000000000010";
    type_cast_1142_wire_constant <= "00000000000000000000000000000001";
    type_cast_1148_wire_constant <= "11111111111111111111111111111111";
    type_cast_1158_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1165_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1176_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1196_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_119_wire_constant <= "0000000000001000";
    type_cast_1206_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1216_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1226_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1236_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1246_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1256_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1290_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_144_wire_constant <= "0000000000001000";
    type_cast_169_wire_constant <= "0000000000001000";
    type_cast_194_wire_constant <= "0000000000001000";
    type_cast_272_wire_constant <= "0000000000001000";
    type_cast_297_wire_constant <= "0000000000001000";
    type_cast_322_wire_constant <= "0000000000001000";
    type_cast_347_wire_constant <= "0000000000001000";
    type_cast_372_wire_constant <= "0000000000001000";
    type_cast_390_wire_constant <= "00000000000000000000000000000011";
    type_cast_406_wire_constant <= "00000000000000000000000000000011";
    type_cast_419_wire_constant <= "00000000000000000000000000000010";
    type_cast_425_wire_constant <= "00000000000000000000000000000001";
    type_cast_431_wire_constant <= "11111111111111111111111111111111";
    type_cast_441_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_448_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_44_wire_constant <= "0000000000001000";
    type_cast_457_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_478_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_496_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_514_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_532_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_550_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_568_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_586_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_608_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_626_wire_constant <= "00000000000000000000000000000010";
    type_cast_632_wire_constant <= "00000000000000000000000000000001";
    type_cast_638_wire_constant <= "11111111111111111111111111111111";
    type_cast_648_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_655_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_666_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_685_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_69_wire_constant <= "0000000000001000";
    type_cast_703_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_721_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_739_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_757_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_775_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_793_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_815_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_857_wire_constant <= "00000000000000000000000000000011";
    type_cast_870_wire_constant <= "00000000000000000000000000000010";
    type_cast_876_wire_constant <= "00000000000000000000000000000001";
    type_cast_882_wire_constant <= "11111111111111111111111111111111";
    type_cast_892_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_899_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_908_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_922_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_927_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_94_wire_constant <= "0000000000001000";
    phi_stmt_1170: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1173_wire & type_cast_1176_wire_constant;
      req <= phi_stmt_1170_req_0 & phi_stmt_1170_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1170",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1170_ack_0,
          idata => idata,
          odata => indvar_1170,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1170
    phi_stmt_453: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_457_wire_constant & type_cast_459_wire;
      req <= phi_stmt_453_req_0 & phi_stmt_453_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_453",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_453_ack_0,
          idata => idata,
          odata => indvar459_453,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_453
    phi_stmt_660: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_663_wire & type_cast_666_wire_constant;
      req <= phi_stmt_660_req_0 & phi_stmt_660_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_660",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_660_ack_0,
          idata => idata,
          odata => indvar443_660,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_660
    phi_stmt_904: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_908_wire_constant & type_cast_910_wire;
      req <= phi_stmt_904_req_0 & phi_stmt_904_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_904",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_904_ack_0,
          idata => idata,
          odata => indvar429_904,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_904
    -- flow-through select operator MUX_1166_inst
    tmp428_1167 <= xx_xop_1160 when (tmp425_1144(0) /=  '0') else type_cast_1165_wire_constant;
    -- flow-through select operator MUX_449_inst
    tmp471_450 <= xx_xop475_443 when (tmp467_427(0) /=  '0') else type_cast_448_wire_constant;
    -- flow-through select operator MUX_656_inst
    tmp457_657 <= xx_xop474_650 when (tmp453_634(0) /=  '0') else type_cast_655_wire_constant;
    -- flow-through select operator MUX_900_inst
    tmp441_901 <= xx_xop473_894 when (tmp437_878(0) /=  '0') else type_cast_899_wire_constant;
    addr_of_1183_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1183_final_reg_req_0;
      addr_of_1183_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1183_final_reg_req_1;
      addr_of_1183_final_reg_ack_1<= rack(0);
      addr_of_1183_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1183_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1182_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx337_1184,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_466_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_466_final_reg_req_0;
      addr_of_466_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_466_final_reg_req_1;
      addr_of_466_final_reg_ack_1<= rack(0);
      addr_of_466_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_466_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_465_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_467,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_673_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_673_final_reg_req_0;
      addr_of_673_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_673_final_reg_req_1;
      addr_of_673_final_reg_ack_1<= rack(0);
      addr_of_673_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_673_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 11,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_672_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx232_674,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_917_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_917_final_reg_req_0;
      addr_of_917_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_917_final_reg_req_1;
      addr_of_917_final_reg_ack_1<= rack(0);
      addr_of_917_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_917_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_916_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx255_918,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_102_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_102_inst_req_0;
      type_cast_102_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_102_inst_req_1;
      type_cast_102_inst_ack_1<= rack(0);
      type_cast_102_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_102_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call19_99,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv20_103,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1115_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1115_inst_req_0;
      type_cast_1115_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1115_inst_req_1;
      type_cast_1115_inst_ack_1<= rack(0);
      type_cast_1115_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1115_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1114_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv321_1116,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_114_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_114_inst_req_0;
      type_cast_114_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_114_inst_req_1;
      type_cast_114_inst_ack_1<= rack(0);
      type_cast_114_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_114_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call23_111,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv26_115,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1153_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1153_inst_req_0;
      type_cast_1153_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1153_inst_req_1;
      type_cast_1153_inst_ack_1<= rack(0);
      type_cast_1153_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1153_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp424x_xop_1150,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_163_1154,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1173_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1173_inst_req_0;
      type_cast_1173_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1173_inst_req_1;
      type_cast_1173_inst_ack_1<= rack(0);
      type_cast_1173_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1173_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1292,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1173_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1191_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1191_inst_req_0;
      type_cast_1191_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1191_inst_req_1;
      type_cast_1191_inst_ack_1<= rack(0);
      type_cast_1191_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1191_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp338_1188,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv341_1192,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1201_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1201_inst_req_0;
      type_cast_1201_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1201_inst_req_1;
      type_cast_1201_inst_ack_1<= rack(0);
      type_cast_1201_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1201_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr344_1198,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv347_1202,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1211_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1211_inst_req_0;
      type_cast_1211_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1211_inst_req_1;
      type_cast_1211_inst_ack_1<= rack(0);
      type_cast_1211_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1211_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr350_1208,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv353_1212,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1221_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1221_inst_req_0;
      type_cast_1221_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1221_inst_req_1;
      type_cast_1221_inst_ack_1<= rack(0);
      type_cast_1221_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1221_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr356_1218,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv359_1222,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1231_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1231_inst_req_0;
      type_cast_1231_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1231_inst_req_1;
      type_cast_1231_inst_ack_1<= rack(0);
      type_cast_1231_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1231_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr362_1228,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv365_1232,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1241_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1241_inst_req_0;
      type_cast_1241_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1241_inst_req_1;
      type_cast_1241_inst_ack_1<= rack(0);
      type_cast_1241_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1241_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr368_1238,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv371_1242,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1251_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1251_inst_req_0;
      type_cast_1251_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1251_inst_req_1;
      type_cast_1251_inst_ack_1<= rack(0);
      type_cast_1251_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1251_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr374_1248,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv377_1252,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1261_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1261_inst_req_0;
      type_cast_1261_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1261_inst_req_1;
      type_cast_1261_inst_ack_1<= rack(0);
      type_cast_1261_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1261_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr380_1258,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv383_1262,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_127_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_127_inst_req_0;
      type_cast_127_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_127_inst_req_1;
      type_cast_127_inst_ack_1<= rack(0);
      type_cast_127_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_127_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call28_124,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_128,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_139_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_139_inst_req_0;
      type_cast_139_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_139_inst_req_1;
      type_cast_139_inst_ack_1<= rack(0);
      type_cast_139_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_139_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call32_136,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv35_140,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_152_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_152_inst_req_0;
      type_cast_152_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_152_inst_req_1;
      type_cast_152_inst_ack_1<= rack(0);
      type_cast_152_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_152_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call37_149,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_153,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_164_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_164_inst_req_0;
      type_cast_164_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_164_inst_req_1;
      type_cast_164_inst_ack_1<= rack(0);
      type_cast_164_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_164_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_161,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_165,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_177_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_177_inst_req_0;
      type_cast_177_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_177_inst_req_1;
      type_cast_177_inst_ack_1<= rack(0);
      type_cast_177_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_177_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_174,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv47_178,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_189_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_189_inst_req_0;
      type_cast_189_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_189_inst_req_1;
      type_cast_189_inst_ack_1<= rack(0);
      type_cast_189_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_189_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call50_186,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv53_190,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_202_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_202_inst_req_0;
      type_cast_202_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_202_inst_req_1;
      type_cast_202_inst_ack_1<= rack(0);
      type_cast_202_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_202_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call55_199,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_203,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_211_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_211_inst_req_0;
      type_cast_211_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_211_inst_req_1;
      type_cast_211_inst_ack_1<= rack(0);
      type_cast_211_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_211_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_58,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv61_212,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_215_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_215_inst_req_0;
      type_cast_215_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_215_inst_req_1;
      type_cast_215_inst_ack_1<= rack(0);
      type_cast_215_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_215_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add12_83,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv63_216,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_219_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_219_inst_req_0;
      type_cast_219_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_219_inst_req_1;
      type_cast_219_inst_ack_1<= rack(0);
      type_cast_219_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_219_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add21_108,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_220,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_233_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_233_inst_req_0;
      type_cast_233_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_233_inst_req_1;
      type_cast_233_inst_ack_1<= rack(0);
      type_cast_233_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_233_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add30_133,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv69_234,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_237_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_237_inst_req_0;
      type_cast_237_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_237_inst_req_1;
      type_cast_237_inst_ack_1<= rack(0);
      type_cast_237_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_237_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add39_158,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv71_238,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_241_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_241_inst_req_0;
      type_cast_241_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_241_inst_req_1;
      type_cast_241_inst_ack_1<= rack(0);
      type_cast_241_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_241_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add48_183,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv74_242,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_245_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_245_inst_req_0;
      type_cast_245_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_245_inst_req_1;
      type_cast_245_inst_ack_1<= rack(0);
      type_cast_245_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_245_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add57_208,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv77_246,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_267_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_267_inst_req_0;
      type_cast_267_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_267_inst_req_1;
      type_cast_267_inst_ack_1<= rack(0);
      type_cast_267_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_267_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call79_264,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv82_268,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_280_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_280_inst_req_0;
      type_cast_280_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_280_inst_req_1;
      type_cast_280_inst_ack_1<= rack(0);
      type_cast_280_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_280_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call84_277,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv85_281,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_292_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_292_inst_req_0;
      type_cast_292_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_292_inst_req_1;
      type_cast_292_inst_ack_1<= rack(0);
      type_cast_292_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_292_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call88_289,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv91_293,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_305_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_305_inst_req_0;
      type_cast_305_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_305_inst_req_1;
      type_cast_305_inst_ack_1<= rack(0);
      type_cast_305_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_305_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call93_302,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv94_306,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_317_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_317_inst_req_0;
      type_cast_317_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_317_inst_req_1;
      type_cast_317_inst_ack_1<= rack(0);
      type_cast_317_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_317_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call97_314,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv100_318,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_330_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_330_inst_req_0;
      type_cast_330_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_330_inst_req_1;
      type_cast_330_inst_ack_1<= rack(0);
      type_cast_330_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_330_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call102_327,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv103_331,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_342_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_342_inst_req_0;
      type_cast_342_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_342_inst_req_1;
      type_cast_342_inst_ack_1<= rack(0);
      type_cast_342_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_342_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call106_339,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv109_343,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_355_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_355_inst_req_0;
      type_cast_355_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_355_inst_req_1;
      type_cast_355_inst_ack_1<= rack(0);
      type_cast_355_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_355_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call111_352,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv112_356,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_367_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_367_inst_req_0;
      type_cast_367_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_367_inst_req_1;
      type_cast_367_inst_ack_1<= rack(0);
      type_cast_367_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_367_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call115_364,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv118_368,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_380_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_380_inst_req_0;
      type_cast_380_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_380_inst_req_1;
      type_cast_380_inst_ack_1<= rack(0);
      type_cast_380_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_380_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call120_377,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv121_381,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_39_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_39_inst_req_0;
      type_cast_39_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_39_inst_req_1;
      type_cast_39_inst_ack_1<= rack(0);
      type_cast_39_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_39_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_36,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1_40,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_436_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_436_inst_req_0;
      type_cast_436_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_436_inst_req_1;
      type_cast_436_inst_ack_1<= rack(0);
      type_cast_436_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_436_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp466x_xop_433,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_25_437,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_459_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_459_inst_req_0;
      type_cast_459_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_459_inst_req_1;
      type_cast_459_inst_ack_1<= rack(0);
      type_cast_459_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_459_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext460_610,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_459_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_473_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_473_inst_req_0;
      type_cast_473_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_473_inst_req_1;
      type_cast_473_inst_ack_1<= rack(0);
      type_cast_473_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_473_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call129_470,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv130_474,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_486_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_486_inst_req_0;
      type_cast_486_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_486_inst_req_1;
      type_cast_486_inst_ack_1<= rack(0);
      type_cast_486_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_486_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call133_483,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv135_487,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_504_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_504_inst_req_0;
      type_cast_504_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_504_inst_req_1;
      type_cast_504_inst_ack_1<= rack(0);
      type_cast_504_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_504_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call139_501,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv141_505,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_522_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_522_inst_req_0;
      type_cast_522_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_522_inst_req_1;
      type_cast_522_inst_ack_1<= rack(0);
      type_cast_522_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_522_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call145_519,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv147_523,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_52_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_52_inst_req_0;
      type_cast_52_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_52_inst_req_1;
      type_cast_52_inst_ack_1<= rack(0);
      type_cast_52_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_52_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_49,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_53,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_540_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_540_inst_req_0;
      type_cast_540_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_540_inst_req_1;
      type_cast_540_inst_ack_1<= rack(0);
      type_cast_540_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_540_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call151_537,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv153_541,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_558_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_558_inst_req_0;
      type_cast_558_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_558_inst_req_1;
      type_cast_558_inst_ack_1<= rack(0);
      type_cast_558_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_558_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call157_555,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv159_559,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_576_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_576_inst_req_0;
      type_cast_576_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_576_inst_req_1;
      type_cast_576_inst_ack_1<= rack(0);
      type_cast_576_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_576_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call163_573,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv165_577,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_594_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_594_inst_req_0;
      type_cast_594_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_594_inst_req_1;
      type_cast_594_inst_ack_1<= rack(0);
      type_cast_594_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_594_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call169_591,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv171_595,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_643_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_643_inst_req_0;
      type_cast_643_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_643_inst_req_1;
      type_cast_643_inst_ack_1<= rack(0);
      type_cast_643_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_643_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp452x_xop_640,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_38_644,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_64_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_64_inst_req_0;
      type_cast_64_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_64_inst_req_1;
      type_cast_64_inst_ack_1<= rack(0);
      type_cast_64_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_64_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_61,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv8_65,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_663_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_663_inst_req_0;
      type_cast_663_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_663_inst_req_1;
      type_cast_663_inst_ack_1<= rack(0);
      type_cast_663_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_663_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext444_817,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_663_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_680_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_680_inst_req_0;
      type_cast_680_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_680_inst_req_1;
      type_cast_680_inst_ack_1<= rack(0);
      type_cast_680_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_680_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call185_677,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv186_681,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_693_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_693_inst_req_0;
      type_cast_693_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_693_inst_req_1;
      type_cast_693_inst_ack_1<= rack(0);
      type_cast_693_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_693_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call189_690,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv191_694,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_711_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_711_inst_req_0;
      type_cast_711_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_711_inst_req_1;
      type_cast_711_inst_ack_1<= rack(0);
      type_cast_711_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_711_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call195_708,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv197_712,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_729_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_729_inst_req_0;
      type_cast_729_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_729_inst_req_1;
      type_cast_729_inst_ack_1<= rack(0);
      type_cast_729_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_729_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call201_726,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv203_730,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_747_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_747_inst_req_0;
      type_cast_747_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_747_inst_req_1;
      type_cast_747_inst_ack_1<= rack(0);
      type_cast_747_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_747_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call207_744,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv209_748,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_765_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_765_inst_req_0;
      type_cast_765_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_765_inst_req_1;
      type_cast_765_inst_ack_1<= rack(0);
      type_cast_765_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_765_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call213_762,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv215_766,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_77_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_77_inst_req_0;
      type_cast_77_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_77_inst_req_1;
      type_cast_77_inst_ack_1<= rack(0);
      type_cast_77_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_77_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call10_74,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv11_78,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_783_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_783_inst_req_0;
      type_cast_783_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_783_inst_req_1;
      type_cast_783_inst_ack_1<= rack(0);
      type_cast_783_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_783_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call219_780,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv221_784,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_801_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_801_inst_req_0;
      type_cast_801_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_801_inst_req_1;
      type_cast_801_inst_ack_1<= rack(0);
      type_cast_801_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_801_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call225_798,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv227_802,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_834_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_834_inst_req_0;
      type_cast_834_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_834_inst_req_1;
      type_cast_834_inst_ack_1<= rack(0);
      type_cast_834_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_834_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add104_336,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv239_835,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_838_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_838_inst_req_0;
      type_cast_838_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_838_inst_req_1;
      type_cast_838_inst_ack_1<= rack(0);
      type_cast_838_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_838_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add113_361,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv241_839,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_842_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_842_inst_req_0;
      type_cast_842_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_842_inst_req_1;
      type_cast_842_inst_ack_1<= rack(0);
      type_cast_842_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_842_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add122_386,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv244_843,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_887_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_887_inst_req_0;
      type_cast_887_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_887_inst_req_1;
      type_cast_887_inst_ack_1<= rack(0);
      type_cast_887_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_887_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp436x_xop_884,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_52_888,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_89_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_89_inst_req_0;
      type_cast_89_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_89_inst_req_1;
      type_cast_89_inst_ack_1<= rack(0);
      type_cast_89_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_89_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call14_86,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_90,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_910_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_910_inst_req_0;
      type_cast_910_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_910_inst_req_1;
      type_cast_910_inst_ack_1<= rack(0);
      type_cast_910_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_910_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext430_929,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_910_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_951_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_951_inst_req_0;
      type_cast_951_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_951_inst_req_1;
      type_cast_951_inst_ack_1<= rack(0);
      type_cast_951_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_951_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_950_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv262_952,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1182_index_1_rename
    process(R_indvar_1181_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_1181_resized;
      ov(13 downto 0) := iv;
      R_indvar_1181_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1182_index_1_resize
    process(indvar_1170) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_1170;
      ov := iv(13 downto 0);
      R_indvar_1181_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1182_root_address_inst
    process(array_obj_ref_1182_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1182_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1182_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_465_index_1_rename
    process(R_indvar459_464_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar459_464_resized;
      ov(13 downto 0) := iv;
      R_indvar459_464_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_465_index_1_resize
    process(indvar459_453) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar459_453;
      ov := iv(13 downto 0);
      R_indvar459_464_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_465_root_address_inst
    process(array_obj_ref_465_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_465_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_465_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_672_index_1_rename
    process(R_indvar443_671_resized) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar443_671_resized;
      ov(10 downto 0) := iv;
      R_indvar443_671_scaled <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_672_index_1_resize
    process(indvar443_660) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar443_660;
      ov := iv(10 downto 0);
      R_indvar443_671_resized <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_672_root_address_inst
    process(array_obj_ref_672_final_offset) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_672_final_offset;
      ov(10 downto 0) := iv;
      array_obj_ref_672_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_916_index_1_rename
    process(R_indvar429_915_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar429_915_resized;
      ov(13 downto 0) := iv;
      R_indvar429_915_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_916_index_1_resize
    process(indvar429_904) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar429_904;
      ov := iv(13 downto 0);
      R_indvar429_915_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_916_root_address_inst
    process(array_obj_ref_916_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_916_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_916_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1187_addr_0
    process(ptr_deref_1187_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1187_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1187_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1187_base_resize
    process(arrayidx337_1184) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx337_1184;
      ov := iv(13 downto 0);
      ptr_deref_1187_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1187_gather_scatter
    process(ptr_deref_1187_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1187_data_0;
      ov(63 downto 0) := iv;
      tmp338_1188 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1187_root_address_inst
    process(ptr_deref_1187_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1187_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1187_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_602_addr_0
    process(ptr_deref_602_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_602_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_602_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_602_base_resize
    process(arrayidx_467) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_467;
      ov := iv(13 downto 0);
      ptr_deref_602_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_602_gather_scatter
    process(add172_600) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add172_600;
      ov(63 downto 0) := iv;
      ptr_deref_602_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_602_root_address_inst
    process(ptr_deref_602_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_602_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_602_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_809_addr_0
    process(ptr_deref_809_root_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_809_root_address;
      ov(10 downto 0) := iv;
      ptr_deref_809_word_address_0 <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_809_base_resize
    process(arrayidx232_674) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx232_674;
      ov := iv(10 downto 0);
      ptr_deref_809_resized_base_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_809_gather_scatter
    process(add228_807) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add228_807;
      ov(63 downto 0) := iv;
      ptr_deref_809_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_809_root_address_inst
    process(ptr_deref_809_resized_base_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_809_resized_base_address;
      ov(10 downto 0) := iv;
      ptr_deref_809_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_920_addr_0
    process(ptr_deref_920_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_920_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_920_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_920_base_resize
    process(arrayidx255_918) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx255_918;
      ov := iv(13 downto 0);
      ptr_deref_920_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_920_gather_scatter
    process(type_cast_922_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_922_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_920_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_920_root_address_inst
    process(ptr_deref_920_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_920_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_920_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1126_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp250409_859;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1126_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1126_branch_req_0,
          ack0 => if_stmt_1126_branch_ack_0,
          ack1 => if_stmt_1126_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1298_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_1297;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1298_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1298_branch_req_0,
          ack0 => if_stmt_1298_branch_ack_0,
          ack1 => if_stmt_1298_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_394_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp417_393;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_394_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_394_branch_req_0,
          ack0 => if_stmt_394_branch_ack_0,
          ack1 => if_stmt_394_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_409_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp180413_408;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_409_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_409_branch_req_0,
          ack0 => if_stmt_409_branch_ack_0,
          ack1 => if_stmt_409_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_616_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond3_615;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_616_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_616_branch_req_0,
          ack0 => if_stmt_616_branch_ack_0,
          ack1 => if_stmt_616_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_823_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond2_822;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_823_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_823_branch_req_0,
          ack0 => if_stmt_823_branch_ack_0,
          ack1 => if_stmt_823_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_860_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp250409_859;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_860_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_860_branch_req_0,
          ack0 => if_stmt_860_branch_ack_0,
          ack1 => if_stmt_860_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_935_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_934;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_935_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_935_branch_req_0,
          ack0 => if_stmt_935_branch_ack_0,
          ack1 => if_stmt_935_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_1149_inst
    process(tmp424_1138) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp424_1138, type_cast_1148_wire_constant, tmp_var);
      tmp424x_xop_1150 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_432_inst
    process(tmp466_421) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp466_421, type_cast_431_wire_constant, tmp_var);
      tmp466x_xop_433 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_639_inst
    process(tmp452_628) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp452_628, type_cast_638_wire_constant, tmp_var);
      tmp452x_xop_640 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_883_inst
    process(tmp436_872) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp436_872, type_cast_882_wire_constant, tmp_var);
      tmp436x_xop_884 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1159_inst
    process(iNsTr_163_1154) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_163_1154, type_cast_1158_wire_constant, tmp_var);
      xx_xop_1160 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1291_inst
    process(indvar_1170) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1170, type_cast_1290_wire_constant, tmp_var);
      indvarx_xnext_1292 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_442_inst
    process(iNsTr_25_437) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_25_437, type_cast_441_wire_constant, tmp_var);
      xx_xop475_443 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_609_inst
    process(indvar459_453) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar459_453, type_cast_608_wire_constant, tmp_var);
      indvarx_xnext460_610 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_649_inst
    process(iNsTr_38_644) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_38_644, type_cast_648_wire_constant, tmp_var);
      xx_xop474_650 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_816_inst
    process(indvar443_660) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar443_660, type_cast_815_wire_constant, tmp_var);
      indvarx_xnext444_817 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_893_inst
    process(iNsTr_52_888) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_52_888, type_cast_892_wire_constant, tmp_var);
      xx_xop473_894 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_928_inst
    process(indvar429_904) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar429_904, type_cast_927_wire_constant, tmp_var);
      indvarx_xnext430_929 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1296_inst
    process(indvarx_xnext_1292, tmp428_1167) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1292, tmp428_1167, tmp_var);
      exitcond1_1297 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_614_inst
    process(indvarx_xnext460_610, tmp471_450) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext460_610, tmp471_450, tmp_var);
      exitcond3_615 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_821_inst
    process(indvarx_xnext444_817, tmp457_657) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext444_817, tmp457_657, tmp_var);
      exitcond2_822 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_933_inst
    process(indvarx_xnext430_929, tmp441_901) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext430_929, tmp441_901, tmp_var);
      exitcond_934 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1137_inst
    process(mul245_853) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul245_853, type_cast_1136_wire_constant, tmp_var);
      tmp424_1138 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_420_inst
    process(mul66_230) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_230, type_cast_419_wire_constant, tmp_var);
      tmp466_421 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_627_inst
    process(mul78_261) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul78_261, type_cast_626_wire_constant, tmp_var);
      tmp452_628 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_871_inst
    process(mul245_853) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul245_853, type_cast_870_wire_constant, tmp_var);
      tmp436_872 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1197_inst
    process(tmp338_1188) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp338_1188, type_cast_1196_wire_constant, tmp_var);
      shr344_1198 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1207_inst
    process(tmp338_1188) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp338_1188, type_cast_1206_wire_constant, tmp_var);
      shr350_1208 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1217_inst
    process(tmp338_1188) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp338_1188, type_cast_1216_wire_constant, tmp_var);
      shr356_1218 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1227_inst
    process(tmp338_1188) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp338_1188, type_cast_1226_wire_constant, tmp_var);
      shr362_1228 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1237_inst
    process(tmp338_1188) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp338_1188, type_cast_1236_wire_constant, tmp_var);
      shr368_1238 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1247_inst
    process(tmp338_1188) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp338_1188, type_cast_1246_wire_constant, tmp_var);
      shr374_1248 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1257_inst
    process(tmp338_1188) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp338_1188, type_cast_1256_wire_constant, tmp_var);
      shr380_1258 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_224_inst
    process(conv63_216, conv61_212) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv63_216, conv61_212, tmp_var);
      mul_225 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_229_inst
    process(mul_225, conv65_220) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_225, conv65_220, tmp_var);
      mul66_230 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_250_inst
    process(conv71_238, conv69_234) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv71_238, conv69_234, tmp_var);
      mul72_251 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_255_inst
    process(mul72_251, conv74_242) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul72_251, conv74_242, tmp_var);
      mul75_256 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_260_inst
    process(mul75_256, conv77_246) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul75_256, conv77_246, tmp_var);
      mul78_261 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_847_inst
    process(conv241_839, conv239_835) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv241_839, conv239_835, tmp_var);
      mul242_848 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_852_inst
    process(mul242_848, conv244_843) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul242_848, conv244_843, tmp_var);
      mul245_853 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_107_inst
    process(shl18_96, conv20_103) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl18_96, conv20_103, tmp_var);
      add21_108 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_132_inst
    process(shl27_121, conv29_128) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl27_121, conv29_128, tmp_var);
      add30_133 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_157_inst
    process(shl36_146, conv38_153) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl36_146, conv38_153, tmp_var);
      add39_158 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_182_inst
    process(shl45_171, conv47_178) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl45_171, conv47_178, tmp_var);
      add48_183 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_207_inst
    process(shl54_196, conv56_203) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl54_196, conv56_203, tmp_var);
      add57_208 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_285_inst
    process(shl83_274, conv85_281) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl83_274, conv85_281, tmp_var);
      add86_286 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_310_inst
    process(shl92_299, conv94_306) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl92_299, conv94_306, tmp_var);
      add95_311 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_335_inst
    process(shl101_324, conv103_331) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl101_324, conv103_331, tmp_var);
      add104_336 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_360_inst
    process(shl110_349, conv112_356) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl110_349, conv112_356, tmp_var);
      add113_361 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_385_inst
    process(shl119_374, conv121_381) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl119_374, conv121_381, tmp_var);
      add122_386 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_57_inst
    process(shl_46, conv3_53) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_46, conv3_53, tmp_var);
      add_58 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_82_inst
    process(shl9_71, conv11_78) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl9_71, conv11_78, tmp_var);
      add12_83 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_491_inst
    process(shl132_480, conv135_487) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl132_480, conv135_487, tmp_var);
      add136_492 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_509_inst
    process(shl138_498, conv141_505) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl138_498, conv141_505, tmp_var);
      add142_510 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_527_inst
    process(shl144_516, conv147_523) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl144_516, conv147_523, tmp_var);
      add148_528 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_545_inst
    process(shl150_534, conv153_541) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl150_534, conv153_541, tmp_var);
      add154_546 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_563_inst
    process(shl156_552, conv159_559) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl156_552, conv159_559, tmp_var);
      add160_564 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_581_inst
    process(shl162_570, conv165_577) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl162_570, conv165_577, tmp_var);
      add166_582 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_599_inst
    process(shl168_588, conv171_595) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl168_588, conv171_595, tmp_var);
      add172_600 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_698_inst
    process(shl188_687, conv191_694) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl188_687, conv191_694, tmp_var);
      add192_699 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_716_inst
    process(shl194_705, conv197_712) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl194_705, conv197_712, tmp_var);
      add198_717 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_734_inst
    process(shl200_723, conv203_730) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl200_723, conv203_730, tmp_var);
      add204_735 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_752_inst
    process(shl206_741, conv209_748) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl206_741, conv209_748, tmp_var);
      add210_753 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_770_inst
    process(shl212_759, conv215_766) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl212_759, conv215_766, tmp_var);
      add216_771 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_788_inst
    process(shl218_777, conv221_784) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl218_777, conv221_784, tmp_var);
      add222_789 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_806_inst
    process(shl224_795, conv227_802) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl224_795, conv227_802, tmp_var);
      add228_807 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_120_inst
    process(conv26_115) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv26_115, type_cast_119_wire_constant, tmp_var);
      shl27_121 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_145_inst
    process(conv35_140) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv35_140, type_cast_144_wire_constant, tmp_var);
      shl36_146 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_170_inst
    process(conv44_165) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv44_165, type_cast_169_wire_constant, tmp_var);
      shl45_171 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_195_inst
    process(conv53_190) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv53_190, type_cast_194_wire_constant, tmp_var);
      shl54_196 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_273_inst
    process(conv82_268) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv82_268, type_cast_272_wire_constant, tmp_var);
      shl83_274 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_298_inst
    process(conv91_293) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv91_293, type_cast_297_wire_constant, tmp_var);
      shl92_299 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_323_inst
    process(conv100_318) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv100_318, type_cast_322_wire_constant, tmp_var);
      shl101_324 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_348_inst
    process(conv109_343) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv109_343, type_cast_347_wire_constant, tmp_var);
      shl110_349 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_373_inst
    process(conv118_368) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv118_368, type_cast_372_wire_constant, tmp_var);
      shl119_374 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_45_inst
    process(conv1_40) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1_40, type_cast_44_wire_constant, tmp_var);
      shl_46 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_70_inst
    process(conv8_65) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv8_65, type_cast_69_wire_constant, tmp_var);
      shl9_71 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_95_inst
    process(conv17_90) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv17_90, type_cast_94_wire_constant, tmp_var);
      shl18_96 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_479_inst
    process(conv130_474) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv130_474, type_cast_478_wire_constant, tmp_var);
      shl132_480 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_497_inst
    process(add136_492) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add136_492, type_cast_496_wire_constant, tmp_var);
      shl138_498 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_515_inst
    process(add142_510) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add142_510, type_cast_514_wire_constant, tmp_var);
      shl144_516 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_533_inst
    process(add148_528) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add148_528, type_cast_532_wire_constant, tmp_var);
      shl150_534 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_551_inst
    process(add154_546) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add154_546, type_cast_550_wire_constant, tmp_var);
      shl156_552 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_569_inst
    process(add160_564) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add160_564, type_cast_568_wire_constant, tmp_var);
      shl162_570 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_587_inst
    process(add166_582) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add166_582, type_cast_586_wire_constant, tmp_var);
      shl168_588 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_686_inst
    process(conv186_681) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv186_681, type_cast_685_wire_constant, tmp_var);
      shl188_687 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_704_inst
    process(add192_699) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add192_699, type_cast_703_wire_constant, tmp_var);
      shl194_705 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_722_inst
    process(add198_717) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add198_717, type_cast_721_wire_constant, tmp_var);
      shl200_723 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_740_inst
    process(add204_735) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add204_735, type_cast_739_wire_constant, tmp_var);
      shl206_741 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_758_inst
    process(add210_753) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add210_753, type_cast_757_wire_constant, tmp_var);
      shl212_759 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_776_inst
    process(add216_771) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add216_771, type_cast_775_wire_constant, tmp_var);
      shl218_777 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_794_inst
    process(add222_789) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add222_789, type_cast_793_wire_constant, tmp_var);
      shl224_795 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_1120_inst
    process(conv321_1116, conv262_952) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv321_1116, conv262_952, tmp_var);
      sub_1121 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1143_inst
    process(tmp424_1138) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp424_1138, type_cast_1142_wire_constant, tmp_var);
      tmp425_1144 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_391_inst
    process(mul66_230) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul66_230, type_cast_390_wire_constant, tmp_var);
      cmp417_393 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_407_inst
    process(mul78_261) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul78_261, type_cast_406_wire_constant, tmp_var);
      cmp180413_408 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_426_inst
    process(tmp466_421) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp466_421, type_cast_425_wire_constant, tmp_var);
      tmp467_427 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_633_inst
    process(tmp452_628) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp452_628, type_cast_632_wire_constant, tmp_var);
      tmp453_634 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_858_inst
    process(mul245_853) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul245_853, type_cast_857_wire_constant, tmp_var);
      cmp250409_859 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_877_inst
    process(tmp436_872) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp436_872, type_cast_876_wire_constant, tmp_var);
      tmp437_878 <= tmp_var; --
    end process;
    -- shared split operator group (94) : array_obj_ref_1182_index_offset 
    ApIntAdd_group_94: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_1181_scaled;
      array_obj_ref_1182_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1182_index_offset_req_0;
      array_obj_ref_1182_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1182_index_offset_req_1;
      array_obj_ref_1182_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_94_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_94_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_94",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 94
    -- shared split operator group (95) : array_obj_ref_465_index_offset 
    ApIntAdd_group_95: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar459_464_scaled;
      array_obj_ref_465_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_465_index_offset_req_0;
      array_obj_ref_465_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_465_index_offset_req_1;
      array_obj_ref_465_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_95_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_95_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_95",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 95
    -- shared split operator group (96) : array_obj_ref_672_index_offset 
    ApIntAdd_group_96: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar443_671_scaled;
      array_obj_ref_672_final_offset <= data_out(10 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_672_index_offset_req_0;
      array_obj_ref_672_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_672_index_offset_req_1;
      array_obj_ref_672_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_96_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_96_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_96",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000100010",
          constant_width => 11,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 96
    -- shared split operator group (97) : array_obj_ref_916_index_offset 
    ApIntAdd_group_97: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar429_915_scaled;
      array_obj_ref_916_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_916_index_offset_req_0;
      array_obj_ref_916_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_916_index_offset_req_1;
      array_obj_ref_916_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_97_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_97_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_97",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 97
    -- unary operator type_cast_1114_inst
    process(call320_1111) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call320_1111, tmp_var);
      type_cast_1114_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_950_inst
    process(call261_946) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call261_946, tmp_var);
      type_cast_950_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_1187_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1187_load_0_req_0;
      ptr_deref_1187_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1187_load_0_req_1;
      ptr_deref_1187_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1187_word_address_0;
      ptr_deref_1187_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(13 downto 0),
          mtag => memory_space_3_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(63 downto 0),
          mtag => memory_space_3_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_602_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_602_store_0_req_0;
      ptr_deref_602_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_602_store_0_req_1;
      ptr_deref_602_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_602_word_address_0;
      data_in <= ptr_deref_602_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_809_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(10 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_809_store_0_req_0;
      ptr_deref_809_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_809_store_0_req_1;
      ptr_deref_809_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_809_word_address_0;
      data_in <= ptr_deref_809_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 11,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(10 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_920_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_920_store_0_req_0;
      ptr_deref_920_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_920_store_0_req_1;
      ptr_deref_920_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_920_word_address_0;
      data_in <= ptr_deref_920_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared inport operator group (0) : RPIPE_Block0_done_1098_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block0_done_1098_inst_req_0;
      RPIPE_Block0_done_1098_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block0_done_1098_inst_req_1;
      RPIPE_Block0_done_1098_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call312_1099 <= data_out(15 downto 0);
      Block0_done_read_0_gI: SplitGuardInterface generic map(name => "Block0_done_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_done_read_0: InputPortRevised -- 
        generic map ( name => "Block0_done_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_done_pipe_read_req(0),
          oack => Block0_done_pipe_read_ack(0),
          odata => Block0_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_Block1_done_1101_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block1_done_1101_inst_req_0;
      RPIPE_Block1_done_1101_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block1_done_1101_inst_req_1;
      RPIPE_Block1_done_1101_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call314_1102 <= data_out(15 downto 0);
      Block1_done_read_1_gI: SplitGuardInterface generic map(name => "Block1_done_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_done_read_1: InputPortRevised -- 
        generic map ( name => "Block1_done_read_1", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_done_pipe_read_req(0),
          oack => Block1_done_pipe_read_ack(0),
          odata => Block1_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_Block2_done_1104_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block2_done_1104_inst_req_0;
      RPIPE_Block2_done_1104_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block2_done_1104_inst_req_1;
      RPIPE_Block2_done_1104_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call316_1105 <= data_out(15 downto 0);
      Block2_done_read_2_gI: SplitGuardInterface generic map(name => "Block2_done_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_done_read_2: InputPortRevised -- 
        generic map ( name => "Block2_done_read_2", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_done_pipe_read_req(0),
          oack => Block2_done_pipe_read_ack(0),
          odata => Block2_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_Block3_done_1107_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block3_done_1107_inst_req_0;
      RPIPE_Block3_done_1107_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block3_done_1107_inst_req_1;
      RPIPE_Block3_done_1107_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call318_1108 <= data_out(15 downto 0);
      Block3_done_read_3_gI: SplitGuardInterface generic map(name => "Block3_done_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_done_read_3: InputPortRevised -- 
        generic map ( name => "Block3_done_read_3", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_done_pipe_read_req(0),
          oack => Block3_done_pipe_read_ack(0),
          odata => Block3_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared inport operator group (4) : RPIPE_ConvTranspose_input_pipe_363_inst RPIPE_ConvTranspose_input_pipe_351_inst RPIPE_ConvTranspose_input_pipe_326_inst RPIPE_ConvTranspose_input_pipe_198_inst RPIPE_ConvTranspose_input_pipe_110_inst RPIPE_ConvTranspose_input_pipe_123_inst RPIPE_ConvTranspose_input_pipe_301_inst RPIPE_ConvTranspose_input_pipe_376_inst RPIPE_ConvTranspose_input_pipe_263_inst RPIPE_ConvTranspose_input_pipe_676_inst RPIPE_ConvTranspose_input_pipe_338_inst RPIPE_ConvTranspose_input_pipe_35_inst RPIPE_ConvTranspose_input_pipe_288_inst RPIPE_ConvTranspose_input_pipe_276_inst RPIPE_ConvTranspose_input_pipe_48_inst RPIPE_ConvTranspose_input_pipe_135_inst RPIPE_ConvTranspose_input_pipe_313_inst RPIPE_ConvTranspose_input_pipe_60_inst RPIPE_ConvTranspose_input_pipe_148_inst RPIPE_ConvTranspose_input_pipe_185_inst RPIPE_ConvTranspose_input_pipe_160_inst RPIPE_ConvTranspose_input_pipe_73_inst RPIPE_ConvTranspose_input_pipe_85_inst RPIPE_ConvTranspose_input_pipe_173_inst RPIPE_ConvTranspose_input_pipe_689_inst RPIPE_ConvTranspose_input_pipe_743_inst RPIPE_ConvTranspose_input_pipe_761_inst RPIPE_ConvTranspose_input_pipe_707_inst RPIPE_ConvTranspose_input_pipe_725_inst RPIPE_ConvTranspose_input_pipe_590_inst RPIPE_ConvTranspose_input_pipe_572_inst RPIPE_ConvTranspose_input_pipe_554_inst RPIPE_ConvTranspose_input_pipe_536_inst RPIPE_ConvTranspose_input_pipe_518_inst RPIPE_ConvTranspose_input_pipe_500_inst RPIPE_ConvTranspose_input_pipe_482_inst RPIPE_ConvTranspose_input_pipe_469_inst RPIPE_ConvTranspose_input_pipe_98_inst RPIPE_ConvTranspose_input_pipe_779_inst RPIPE_ConvTranspose_input_pipe_797_inst 
    InportGroup_4: Block -- 
      signal data_out: std_logic_vector(319 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 39 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 39 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 39 downto 0);
      signal guard_vector : std_logic_vector( 39 downto 0);
      constant outBUFs : IntegerArray(39 downto 0) := (39 => 1, 38 => 1, 37 => 1, 36 => 1, 35 => 1, 34 => 1, 33 => 1, 32 => 1, 31 => 1, 30 => 1, 29 => 1, 28 => 1, 27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(39 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false, 28 => false, 29 => false, 30 => false, 31 => false, 32 => false, 33 => false, 34 => false, 35 => false, 36 => false, 37 => false, 38 => false, 39 => false);
      constant guardBuffering: IntegerArray(39 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2, 28 => 2, 29 => 2, 30 => 2, 31 => 2, 32 => 2, 33 => 2, 34 => 2, 35 => 2, 36 => 2, 37 => 2, 38 => 2, 39 => 2);
      -- 
    begin -- 
      reqL_unguarded(39) <= RPIPE_ConvTranspose_input_pipe_363_inst_req_0;
      reqL_unguarded(38) <= RPIPE_ConvTranspose_input_pipe_351_inst_req_0;
      reqL_unguarded(37) <= RPIPE_ConvTranspose_input_pipe_326_inst_req_0;
      reqL_unguarded(36) <= RPIPE_ConvTranspose_input_pipe_198_inst_req_0;
      reqL_unguarded(35) <= RPIPE_ConvTranspose_input_pipe_110_inst_req_0;
      reqL_unguarded(34) <= RPIPE_ConvTranspose_input_pipe_123_inst_req_0;
      reqL_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_301_inst_req_0;
      reqL_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_376_inst_req_0;
      reqL_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_263_inst_req_0;
      reqL_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_676_inst_req_0;
      reqL_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_338_inst_req_0;
      reqL_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_35_inst_req_0;
      reqL_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_288_inst_req_0;
      reqL_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_276_inst_req_0;
      reqL_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_48_inst_req_0;
      reqL_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_135_inst_req_0;
      reqL_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_313_inst_req_0;
      reqL_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_60_inst_req_0;
      reqL_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_148_inst_req_0;
      reqL_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_185_inst_req_0;
      reqL_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_160_inst_req_0;
      reqL_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_73_inst_req_0;
      reqL_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_85_inst_req_0;
      reqL_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_173_inst_req_0;
      reqL_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_689_inst_req_0;
      reqL_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_743_inst_req_0;
      reqL_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_761_inst_req_0;
      reqL_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_707_inst_req_0;
      reqL_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_725_inst_req_0;
      reqL_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_590_inst_req_0;
      reqL_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_572_inst_req_0;
      reqL_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_554_inst_req_0;
      reqL_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_536_inst_req_0;
      reqL_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_518_inst_req_0;
      reqL_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_500_inst_req_0;
      reqL_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_482_inst_req_0;
      reqL_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_469_inst_req_0;
      reqL_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_98_inst_req_0;
      reqL_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_779_inst_req_0;
      reqL_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_797_inst_req_0;
      RPIPE_ConvTranspose_input_pipe_363_inst_ack_0 <= ackL_unguarded(39);
      RPIPE_ConvTranspose_input_pipe_351_inst_ack_0 <= ackL_unguarded(38);
      RPIPE_ConvTranspose_input_pipe_326_inst_ack_0 <= ackL_unguarded(37);
      RPIPE_ConvTranspose_input_pipe_198_inst_ack_0 <= ackL_unguarded(36);
      RPIPE_ConvTranspose_input_pipe_110_inst_ack_0 <= ackL_unguarded(35);
      RPIPE_ConvTranspose_input_pipe_123_inst_ack_0 <= ackL_unguarded(34);
      RPIPE_ConvTranspose_input_pipe_301_inst_ack_0 <= ackL_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_376_inst_ack_0 <= ackL_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_263_inst_ack_0 <= ackL_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_676_inst_ack_0 <= ackL_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_338_inst_ack_0 <= ackL_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_35_inst_ack_0 <= ackL_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_288_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_276_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_48_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_135_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_313_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_60_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_148_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_185_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_160_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_73_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_85_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_173_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_689_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_743_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_761_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_707_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_725_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_590_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_572_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_554_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_536_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_518_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_500_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_482_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_469_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_98_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_779_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_797_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(39) <= RPIPE_ConvTranspose_input_pipe_363_inst_req_1;
      reqR_unguarded(38) <= RPIPE_ConvTranspose_input_pipe_351_inst_req_1;
      reqR_unguarded(37) <= RPIPE_ConvTranspose_input_pipe_326_inst_req_1;
      reqR_unguarded(36) <= RPIPE_ConvTranspose_input_pipe_198_inst_req_1;
      reqR_unguarded(35) <= RPIPE_ConvTranspose_input_pipe_110_inst_req_1;
      reqR_unguarded(34) <= RPIPE_ConvTranspose_input_pipe_123_inst_req_1;
      reqR_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_301_inst_req_1;
      reqR_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_376_inst_req_1;
      reqR_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_263_inst_req_1;
      reqR_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_676_inst_req_1;
      reqR_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_338_inst_req_1;
      reqR_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_35_inst_req_1;
      reqR_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_288_inst_req_1;
      reqR_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_276_inst_req_1;
      reqR_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_48_inst_req_1;
      reqR_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_135_inst_req_1;
      reqR_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_313_inst_req_1;
      reqR_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_60_inst_req_1;
      reqR_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_148_inst_req_1;
      reqR_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_185_inst_req_1;
      reqR_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_160_inst_req_1;
      reqR_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_73_inst_req_1;
      reqR_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_85_inst_req_1;
      reqR_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_173_inst_req_1;
      reqR_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_689_inst_req_1;
      reqR_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_743_inst_req_1;
      reqR_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_761_inst_req_1;
      reqR_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_707_inst_req_1;
      reqR_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_725_inst_req_1;
      reqR_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_590_inst_req_1;
      reqR_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_572_inst_req_1;
      reqR_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_554_inst_req_1;
      reqR_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_536_inst_req_1;
      reqR_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_518_inst_req_1;
      reqR_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_500_inst_req_1;
      reqR_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_482_inst_req_1;
      reqR_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_469_inst_req_1;
      reqR_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_98_inst_req_1;
      reqR_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_779_inst_req_1;
      reqR_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_797_inst_req_1;
      RPIPE_ConvTranspose_input_pipe_363_inst_ack_1 <= ackR_unguarded(39);
      RPIPE_ConvTranspose_input_pipe_351_inst_ack_1 <= ackR_unguarded(38);
      RPIPE_ConvTranspose_input_pipe_326_inst_ack_1 <= ackR_unguarded(37);
      RPIPE_ConvTranspose_input_pipe_198_inst_ack_1 <= ackR_unguarded(36);
      RPIPE_ConvTranspose_input_pipe_110_inst_ack_1 <= ackR_unguarded(35);
      RPIPE_ConvTranspose_input_pipe_123_inst_ack_1 <= ackR_unguarded(34);
      RPIPE_ConvTranspose_input_pipe_301_inst_ack_1 <= ackR_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_376_inst_ack_1 <= ackR_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_263_inst_ack_1 <= ackR_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_676_inst_ack_1 <= ackR_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_338_inst_ack_1 <= ackR_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_35_inst_ack_1 <= ackR_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_288_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_276_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_48_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_135_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_313_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_60_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_148_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_185_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_160_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_73_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_85_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_173_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_689_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_743_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_761_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_707_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_725_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_590_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_572_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_554_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_536_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_518_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_500_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_482_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_469_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_98_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_779_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_797_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      guard_vector(34)  <=  '1';
      guard_vector(35)  <=  '1';
      guard_vector(36)  <=  '1';
      guard_vector(37)  <=  '1';
      guard_vector(38)  <=  '1';
      guard_vector(39)  <=  '1';
      call115_364 <= data_out(319 downto 312);
      call111_352 <= data_out(311 downto 304);
      call102_327 <= data_out(303 downto 296);
      call55_199 <= data_out(295 downto 288);
      call23_111 <= data_out(287 downto 280);
      call28_124 <= data_out(279 downto 272);
      call93_302 <= data_out(271 downto 264);
      call120_377 <= data_out(263 downto 256);
      call79_264 <= data_out(255 downto 248);
      call185_677 <= data_out(247 downto 240);
      call106_339 <= data_out(239 downto 232);
      call_36 <= data_out(231 downto 224);
      call88_289 <= data_out(223 downto 216);
      call84_277 <= data_out(215 downto 208);
      call2_49 <= data_out(207 downto 200);
      call32_136 <= data_out(199 downto 192);
      call97_314 <= data_out(191 downto 184);
      call5_61 <= data_out(183 downto 176);
      call37_149 <= data_out(175 downto 168);
      call50_186 <= data_out(167 downto 160);
      call41_161 <= data_out(159 downto 152);
      call10_74 <= data_out(151 downto 144);
      call14_86 <= data_out(143 downto 136);
      call46_174 <= data_out(135 downto 128);
      call189_690 <= data_out(127 downto 120);
      call207_744 <= data_out(119 downto 112);
      call213_762 <= data_out(111 downto 104);
      call195_708 <= data_out(103 downto 96);
      call201_726 <= data_out(95 downto 88);
      call169_591 <= data_out(87 downto 80);
      call163_573 <= data_out(79 downto 72);
      call157_555 <= data_out(71 downto 64);
      call151_537 <= data_out(63 downto 56);
      call145_519 <= data_out(55 downto 48);
      call139_501 <= data_out(47 downto 40);
      call133_483 <= data_out(39 downto 32);
      call129_470 <= data_out(31 downto 24);
      call19_99 <= data_out(23 downto 16);
      call219_780 <= data_out(15 downto 8);
      call225_798 <= data_out(7 downto 0);
      ConvTranspose_input_pipe_read_4_gI: SplitGuardInterface generic map(name => "ConvTranspose_input_pipe_read_4_gI", nreqs => 40, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_input_pipe_read_4: InputPortRevised -- 
        generic map ( name => "ConvTranspose_input_pipe_read_4", data_width => 8,  num_reqs => 40,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => ConvTranspose_input_pipe_pipe_read_req(0),
          oack => ConvTranspose_input_pipe_pipe_read_ack(0),
          odata => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 4
    -- shared outport operator group (0) : WPIPE_Block0_start_953_inst WPIPE_Block0_start_956_inst WPIPE_Block0_start_959_inst WPIPE_Block0_start_962_inst WPIPE_Block0_start_965_inst WPIPE_Block0_start_968_inst WPIPE_Block0_start_971_inst WPIPE_Block0_start_974_inst WPIPE_Block0_start_977_inst WPIPE_Block0_start_980_inst WPIPE_Block0_start_983_inst WPIPE_Block0_start_986_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(191 downto 0);
      signal sample_req, sample_ack : BooleanArray( 11 downto 0);
      signal update_req, update_ack : BooleanArray( 11 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 11 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 11 downto 0);
      signal guard_vector : std_logic_vector( 11 downto 0);
      constant inBUFs : IntegerArray(11 downto 0) := (11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(11 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false);
      constant guardBuffering: IntegerArray(11 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2);
      -- 
    begin -- 
      sample_req_unguarded(11) <= WPIPE_Block0_start_953_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block0_start_956_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block0_start_959_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block0_start_962_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block0_start_965_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block0_start_968_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block0_start_971_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block0_start_974_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block0_start_977_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block0_start_980_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block0_start_983_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block0_start_986_inst_req_0;
      WPIPE_Block0_start_953_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block0_start_956_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block0_start_959_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block0_start_962_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block0_start_965_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block0_start_968_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block0_start_971_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block0_start_974_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block0_start_977_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block0_start_980_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block0_start_983_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block0_start_986_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(11) <= WPIPE_Block0_start_953_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block0_start_956_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block0_start_959_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block0_start_962_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block0_start_965_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block0_start_968_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block0_start_971_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block0_start_974_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block0_start_977_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block0_start_980_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block0_start_983_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block0_start_986_inst_req_1;
      WPIPE_Block0_start_953_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block0_start_956_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block0_start_959_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block0_start_962_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block0_start_965_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block0_start_968_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block0_start_971_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block0_start_974_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block0_start_977_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block0_start_980_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block0_start_983_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block0_start_986_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      data_in <= add_58 & add12_83 & add21_108 & add30_133 & add39_158 & add48_183 & add57_208 & add86_286 & add95_311 & add104_336 & add113_361 & add122_386;
      Block0_start_write_0_gI: SplitGuardInterface generic map(name => "Block0_start_write_0_gI", nreqs => 12, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_start_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_start", data_width => 16, num_reqs => 12, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_start_pipe_write_req(0),
          oack => Block0_start_pipe_write_ack(0),
          odata => Block0_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_Block1_start_989_inst WPIPE_Block1_start_992_inst WPIPE_Block1_start_995_inst WPIPE_Block1_start_998_inst WPIPE_Block1_start_1001_inst WPIPE_Block1_start_1004_inst WPIPE_Block1_start_1007_inst WPIPE_Block1_start_1010_inst WPIPE_Block1_start_1013_inst WPIPE_Block1_start_1016_inst WPIPE_Block1_start_1019_inst WPIPE_Block1_start_1022_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(191 downto 0);
      signal sample_req, sample_ack : BooleanArray( 11 downto 0);
      signal update_req, update_ack : BooleanArray( 11 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 11 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 11 downto 0);
      signal guard_vector : std_logic_vector( 11 downto 0);
      constant inBUFs : IntegerArray(11 downto 0) := (11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(11 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false);
      constant guardBuffering: IntegerArray(11 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2);
      -- 
    begin -- 
      sample_req_unguarded(11) <= WPIPE_Block1_start_989_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block1_start_992_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block1_start_995_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block1_start_998_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block1_start_1001_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block1_start_1004_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block1_start_1007_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block1_start_1010_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block1_start_1013_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block1_start_1016_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block1_start_1019_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block1_start_1022_inst_req_0;
      WPIPE_Block1_start_989_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block1_start_992_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block1_start_995_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block1_start_998_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block1_start_1001_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block1_start_1004_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block1_start_1007_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block1_start_1010_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block1_start_1013_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block1_start_1016_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block1_start_1019_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block1_start_1022_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(11) <= WPIPE_Block1_start_989_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block1_start_992_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block1_start_995_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block1_start_998_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block1_start_1001_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block1_start_1004_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block1_start_1007_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block1_start_1010_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block1_start_1013_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block1_start_1016_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block1_start_1019_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block1_start_1022_inst_req_1;
      WPIPE_Block1_start_989_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block1_start_992_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block1_start_995_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block1_start_998_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block1_start_1001_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block1_start_1004_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block1_start_1007_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block1_start_1010_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block1_start_1013_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block1_start_1016_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block1_start_1019_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block1_start_1022_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      data_in <= add_58 & add12_83 & add21_108 & add30_133 & add39_158 & add48_183 & add57_208 & add86_286 & add95_311 & add104_336 & add113_361 & add122_386;
      Block1_start_write_1_gI: SplitGuardInterface generic map(name => "Block1_start_write_1_gI", nreqs => 12, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_start_write_1: OutputPortRevised -- 
        generic map ( name => "Block1_start", data_width => 16, num_reqs => 12, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_start_pipe_write_req(0),
          oack => Block1_start_pipe_write_ack(0),
          odata => Block1_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_Block2_start_1025_inst WPIPE_Block2_start_1028_inst WPIPE_Block2_start_1031_inst WPIPE_Block2_start_1034_inst WPIPE_Block2_start_1037_inst WPIPE_Block2_start_1040_inst WPIPE_Block2_start_1043_inst WPIPE_Block2_start_1046_inst WPIPE_Block2_start_1049_inst WPIPE_Block2_start_1052_inst WPIPE_Block2_start_1055_inst WPIPE_Block2_start_1058_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(191 downto 0);
      signal sample_req, sample_ack : BooleanArray( 11 downto 0);
      signal update_req, update_ack : BooleanArray( 11 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 11 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 11 downto 0);
      signal guard_vector : std_logic_vector( 11 downto 0);
      constant inBUFs : IntegerArray(11 downto 0) := (11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(11 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false);
      constant guardBuffering: IntegerArray(11 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2);
      -- 
    begin -- 
      sample_req_unguarded(11) <= WPIPE_Block2_start_1025_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block2_start_1028_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block2_start_1031_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block2_start_1034_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block2_start_1037_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block2_start_1040_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block2_start_1043_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block2_start_1046_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block2_start_1049_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block2_start_1052_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block2_start_1055_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block2_start_1058_inst_req_0;
      WPIPE_Block2_start_1025_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block2_start_1028_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block2_start_1031_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block2_start_1034_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block2_start_1037_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block2_start_1040_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block2_start_1043_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block2_start_1046_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block2_start_1049_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block2_start_1052_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block2_start_1055_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block2_start_1058_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(11) <= WPIPE_Block2_start_1025_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block2_start_1028_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block2_start_1031_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block2_start_1034_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block2_start_1037_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block2_start_1040_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block2_start_1043_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block2_start_1046_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block2_start_1049_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block2_start_1052_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block2_start_1055_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block2_start_1058_inst_req_1;
      WPIPE_Block2_start_1025_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block2_start_1028_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block2_start_1031_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block2_start_1034_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block2_start_1037_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block2_start_1040_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block2_start_1043_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block2_start_1046_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block2_start_1049_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block2_start_1052_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block2_start_1055_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block2_start_1058_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      data_in <= add_58 & add12_83 & add21_108 & add30_133 & add39_158 & add48_183 & add57_208 & add86_286 & add95_311 & add104_336 & add113_361 & add122_386;
      Block2_start_write_2_gI: SplitGuardInterface generic map(name => "Block2_start_write_2_gI", nreqs => 12, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_start_write_2: OutputPortRevised -- 
        generic map ( name => "Block2_start", data_width => 16, num_reqs => 12, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_start_pipe_write_req(0),
          oack => Block2_start_pipe_write_ack(0),
          odata => Block2_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_Block3_start_1061_inst WPIPE_Block3_start_1064_inst WPIPE_Block3_start_1067_inst WPIPE_Block3_start_1070_inst WPIPE_Block3_start_1073_inst WPIPE_Block3_start_1076_inst WPIPE_Block3_start_1079_inst WPIPE_Block3_start_1082_inst WPIPE_Block3_start_1085_inst WPIPE_Block3_start_1088_inst WPIPE_Block3_start_1091_inst WPIPE_Block3_start_1094_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(191 downto 0);
      signal sample_req, sample_ack : BooleanArray( 11 downto 0);
      signal update_req, update_ack : BooleanArray( 11 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 11 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 11 downto 0);
      signal guard_vector : std_logic_vector( 11 downto 0);
      constant inBUFs : IntegerArray(11 downto 0) := (11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(11 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false);
      constant guardBuffering: IntegerArray(11 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2);
      -- 
    begin -- 
      sample_req_unguarded(11) <= WPIPE_Block3_start_1061_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block3_start_1064_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block3_start_1067_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block3_start_1070_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block3_start_1073_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block3_start_1076_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block3_start_1079_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block3_start_1082_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block3_start_1085_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block3_start_1088_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block3_start_1091_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block3_start_1094_inst_req_0;
      WPIPE_Block3_start_1061_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block3_start_1064_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block3_start_1067_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block3_start_1070_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block3_start_1073_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block3_start_1076_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block3_start_1079_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block3_start_1082_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block3_start_1085_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block3_start_1088_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block3_start_1091_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block3_start_1094_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(11) <= WPIPE_Block3_start_1061_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block3_start_1064_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block3_start_1067_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block3_start_1070_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block3_start_1073_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block3_start_1076_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block3_start_1079_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block3_start_1082_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block3_start_1085_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block3_start_1088_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block3_start_1091_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block3_start_1094_inst_req_1;
      WPIPE_Block3_start_1061_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block3_start_1064_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block3_start_1067_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block3_start_1070_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block3_start_1073_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block3_start_1076_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block3_start_1079_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block3_start_1082_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block3_start_1085_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block3_start_1088_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block3_start_1091_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block3_start_1094_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      data_in <= add_58 & add12_83 & add21_108 & add30_133 & add39_158 & add48_183 & add57_208 & add86_286 & add95_311 & add104_336 & add113_361 & add122_386;
      Block3_start_write_3_gI: SplitGuardInterface generic map(name => "Block3_start_write_3_gI", nreqs => 12, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_start_write_3: OutputPortRevised -- 
        generic map ( name => "Block3_start", data_width => 16, num_reqs => 12, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_start_pipe_write_req(0),
          oack => Block3_start_pipe_write_ack(0),
          odata => Block3_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared outport operator group (4) : WPIPE_ConvTranspose_output_pipe_1269_inst WPIPE_ConvTranspose_output_pipe_1263_inst WPIPE_ConvTranspose_output_pipe_1266_inst WPIPE_ConvTranspose_output_pipe_1284_inst WPIPE_ConvTranspose_output_pipe_1281_inst WPIPE_ConvTranspose_output_pipe_1278_inst WPIPE_ConvTranspose_output_pipe_1275_inst WPIPE_ConvTranspose_output_pipe_1272_inst 
    OutportGroup_4: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 7 downto 0);
      signal update_req, update_ack : BooleanArray( 7 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 7 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      sample_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1269_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1263_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1266_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1284_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1281_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1278_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1275_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1272_inst_req_0;
      WPIPE_ConvTranspose_output_pipe_1269_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1263_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1266_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1284_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1281_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1278_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1275_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1272_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1269_inst_req_1;
      update_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1263_inst_req_1;
      update_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1266_inst_req_1;
      update_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1284_inst_req_1;
      update_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1281_inst_req_1;
      update_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1278_inst_req_1;
      update_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1275_inst_req_1;
      update_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1272_inst_req_1;
      WPIPE_ConvTranspose_output_pipe_1269_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1263_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1266_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1284_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1281_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1278_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1275_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1272_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      data_in <= conv371_1242 & conv383_1262 & conv377_1252 & conv341_1192 & conv347_1202 & conv353_1212 & conv359_1222 & conv365_1232;
      ConvTranspose_output_pipe_write_4_gI: SplitGuardInterface generic map(name => "ConvTranspose_output_pipe_write_4_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_output_pipe_write_4: OutputPortRevised -- 
        generic map ( name => "ConvTranspose_output_pipe", data_width => 8, num_reqs => 8, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => ConvTranspose_output_pipe_pipe_write_req(0),
          oack => ConvTranspose_output_pipe_pipe_write_ack(0),
          odata => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 4
    -- shared outport operator group (5) : WPIPE_elapsed_time_pipe_1122_inst 
    OutportGroup_5: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1122_inst_req_0;
      WPIPE_elapsed_time_pipe_1122_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1122_inst_req_1;
      WPIPE_elapsed_time_pipe_1122_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= sub_1121;
      elapsed_time_pipe_write_5_gI: SplitGuardInterface generic map(name => "elapsed_time_pipe_write_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      elapsed_time_pipe_write_5: OutputPortRevised -- 
        generic map ( name => "elapsed_time_pipe", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => elapsed_time_pipe_pipe_write_req(0),
          oack => elapsed_time_pipe_pipe_write_ack(0),
          odata => elapsed_time_pipe_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 5
    -- shared call operator group (0) : call_stmt_946_call call_stmt_1111_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_946_call_req_0;
      reqL_unguarded(0) <= call_stmt_1111_call_req_0;
      call_stmt_946_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1111_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_946_call_req_1;
      reqR_unguarded(0) <= call_stmt_1111_call_req_1;
      call_stmt_946_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1111_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call261_946 <= data_out(127 downto 64);
      call320_1111 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end convTranspose_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeA is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeA;
architecture convTransposeA_arch of convTransposeA is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeA_CP_3352_start: Boolean;
  signal convTransposeA_CP_3352_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block0_start_1326_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1317_inst_ack_1 : boolean;
  signal phi_stmt_1405_ack_0 : boolean;
  signal RPIPE_Block0_start_1314_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1323_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1326_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1317_inst_ack_0 : boolean;
  signal type_cast_1618_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1317_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1320_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1329_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1329_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1320_inst_req_1 : boolean;
  signal type_cast_1601_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1326_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1314_inst_ack_1 : boolean;
  signal type_cast_1411_inst_req_1 : boolean;
  signal type_cast_1411_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1320_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1317_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1314_inst_req_1 : boolean;
  signal phi_stmt_1405_req_1 : boolean;
  signal RPIPE_Block0_start_1323_inst_req_0 : boolean;
  signal type_cast_1471_inst_req_0 : boolean;
  signal phi_stmt_1405_req_0 : boolean;
  signal RPIPE_Block0_start_1323_inst_ack_1 : boolean;
  signal if_stmt_1625_branch_req_0 : boolean;
  signal type_cast_1601_inst_req_0 : boolean;
  signal phi_stmt_1398_ack_0 : boolean;
  signal type_cast_1601_inst_ack_1 : boolean;
  signal type_cast_1601_inst_req_1 : boolean;
  signal if_stmt_1625_branch_ack_1 : boolean;
  signal if_stmt_1625_branch_ack_0 : boolean;
  signal type_cast_1471_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1314_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1323_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1326_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1320_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1329_inst_req_1 : boolean;
  signal phi_stmt_1398_req_0 : boolean;
  signal type_cast_1618_inst_req_0 : boolean;
  signal type_cast_1618_inst_ack_0 : boolean;
  signal type_cast_1471_inst_req_1 : boolean;
  signal type_cast_1471_inst_ack_1 : boolean;
  signal type_cast_1618_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1329_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1332_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1332_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1332_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1332_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1335_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1335_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1335_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1335_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1338_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1338_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1338_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1338_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1341_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1341_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1341_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1341_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1344_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1344_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1344_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1344_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1347_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1347_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1347_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1347_inst_ack_1 : boolean;
  signal type_cast_1352_inst_req_0 : boolean;
  signal type_cast_1352_inst_ack_0 : boolean;
  signal type_cast_1352_inst_req_1 : boolean;
  signal type_cast_1352_inst_ack_1 : boolean;
  signal type_cast_1356_inst_req_0 : boolean;
  signal type_cast_1356_inst_ack_0 : boolean;
  signal type_cast_1356_inst_req_1 : boolean;
  signal type_cast_1356_inst_ack_1 : boolean;
  signal type_cast_1366_inst_req_0 : boolean;
  signal type_cast_1366_inst_ack_0 : boolean;
  signal type_cast_1366_inst_req_1 : boolean;
  signal type_cast_1366_inst_ack_1 : boolean;
  signal type_cast_1411_inst_ack_0 : boolean;
  signal type_cast_1493_inst_req_0 : boolean;
  signal phi_stmt_1465_ack_0 : boolean;
  signal type_cast_1493_inst_ack_0 : boolean;
  signal type_cast_1493_inst_req_1 : boolean;
  signal type_cast_1493_inst_ack_1 : boolean;
  signal type_cast_1411_inst_req_0 : boolean;
  signal type_cast_1507_inst_req_0 : boolean;
  signal type_cast_1507_inst_ack_0 : boolean;
  signal type_cast_1592_inst_ack_1 : boolean;
  signal type_cast_1507_inst_req_1 : boolean;
  signal phi_stmt_1465_req_0 : boolean;
  signal type_cast_1507_inst_ack_1 : boolean;
  signal WPIPE_Block0_done_1633_inst_ack_1 : boolean;
  signal WPIPE_Block0_done_1633_inst_req_1 : boolean;
  signal type_cast_1592_inst_req_1 : boolean;
  signal phi_stmt_1398_req_1 : boolean;
  signal type_cast_1404_inst_ack_1 : boolean;
  signal type_cast_1404_inst_req_1 : boolean;
  signal array_obj_ref_1513_index_offset_req_0 : boolean;
  signal array_obj_ref_1513_index_offset_ack_0 : boolean;
  signal array_obj_ref_1513_index_offset_req_1 : boolean;
  signal array_obj_ref_1513_index_offset_ack_1 : boolean;
  signal addr_of_1514_final_reg_req_0 : boolean;
  signal addr_of_1514_final_reg_ack_0 : boolean;
  signal addr_of_1514_final_reg_req_1 : boolean;
  signal addr_of_1514_final_reg_ack_1 : boolean;
  signal WPIPE_Block0_done_1633_inst_ack_0 : boolean;
  signal WPIPE_Block0_done_1633_inst_req_0 : boolean;
  signal type_cast_1404_inst_ack_0 : boolean;
  signal type_cast_1404_inst_req_0 : boolean;
  signal phi_stmt_1465_req_1 : boolean;
  signal ptr_deref_1518_load_0_req_0 : boolean;
  signal ptr_deref_1518_load_0_ack_0 : boolean;
  signal ptr_deref_1518_load_0_req_1 : boolean;
  signal ptr_deref_1518_load_0_ack_1 : boolean;
  signal type_cast_1523_inst_req_0 : boolean;
  signal type_cast_1523_inst_ack_0 : boolean;
  signal type_cast_1523_inst_req_1 : boolean;
  signal type_cast_1523_inst_ack_1 : boolean;
  signal type_cast_1537_inst_req_0 : boolean;
  signal type_cast_1537_inst_ack_0 : boolean;
  signal type_cast_1537_inst_req_1 : boolean;
  signal type_cast_1537_inst_ack_1 : boolean;
  signal array_obj_ref_1543_index_offset_req_0 : boolean;
  signal array_obj_ref_1543_index_offset_ack_0 : boolean;
  signal array_obj_ref_1543_index_offset_req_1 : boolean;
  signal array_obj_ref_1543_index_offset_ack_1 : boolean;
  signal addr_of_1544_final_reg_req_0 : boolean;
  signal addr_of_1544_final_reg_ack_0 : boolean;
  signal addr_of_1544_final_reg_req_1 : boolean;
  signal addr_of_1544_final_reg_ack_1 : boolean;
  signal ptr_deref_1547_store_0_req_0 : boolean;
  signal ptr_deref_1547_store_0_ack_0 : boolean;
  signal ptr_deref_1547_store_0_req_1 : boolean;
  signal ptr_deref_1547_store_0_ack_1 : boolean;
  signal type_cast_1553_inst_req_0 : boolean;
  signal type_cast_1553_inst_ack_0 : boolean;
  signal type_cast_1553_inst_req_1 : boolean;
  signal type_cast_1553_inst_ack_1 : boolean;
  signal if_stmt_1568_branch_req_0 : boolean;
  signal if_stmt_1568_branch_ack_1 : boolean;
  signal if_stmt_1568_branch_ack_0 : boolean;
  signal type_cast_1592_inst_req_0 : boolean;
  signal type_cast_1592_inst_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeA_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeA_CP_3352_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeA_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_3352_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeA_CP_3352_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_3352_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeA_CP_3352: Block -- control-path 
    signal convTransposeA_CP_3352_elements: BooleanArray(87 downto 0);
    -- 
  begin -- 
    convTransposeA_CP_3352_elements(0) <= convTransposeA_CP_3352_start;
    convTransposeA_CP_3352_symbol <= convTransposeA_CP_3352_elements(67);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1314_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1312/$entry
      -- CP-element group 0: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/$entry
      -- CP-element group 0: 	 branch_block_stmt_1312/branch_block_stmt_1312__entry__
      -- CP-element group 0: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348__entry__
      -- CP-element group 0: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1314_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1314_Sample/rr
      -- CP-element group 0: 	 $entry
      -- 
    rr_3400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(0), ack => RPIPE_Block0_start_1314_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1314_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1314_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1314_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1314_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1314_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1314_update_start_
      -- 
    ra_3401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1314_inst_ack_0, ack => convTransposeA_CP_3352_elements(1)); -- 
    cr_3405_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3405_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(1), ack => RPIPE_Block0_start_1314_inst_req_1); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1317_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1314_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1317_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1317_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1314_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1314_Update/$exit
      -- 
    ca_3406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1314_inst_ack_1, ack => convTransposeA_CP_3352_elements(2)); -- 
    rr_3414_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3414_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(2), ack => RPIPE_Block0_start_1317_inst_req_0); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1317_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1317_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1317_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1317_Update/cr
      -- CP-element group 3: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1317_update_start_
      -- CP-element group 3: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1317_Update/$entry
      -- 
    ra_3415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1317_inst_ack_0, ack => convTransposeA_CP_3352_elements(3)); -- 
    cr_3419_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3419_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(3), ack => RPIPE_Block0_start_1317_inst_req_1); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1320_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1317_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1317_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1320_Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1317_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1320_sample_start_
      -- 
    ca_3420_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1317_inst_ack_1, ack => convTransposeA_CP_3352_elements(4)); -- 
    rr_3428_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3428_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(4), ack => RPIPE_Block0_start_1320_inst_req_0); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1320_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1320_update_start_
      -- CP-element group 5: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1320_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1320_Update/cr
      -- CP-element group 5: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1320_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1320_Sample/ra
      -- 
    ra_3429_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1320_inst_ack_0, ack => convTransposeA_CP_3352_elements(5)); -- 
    cr_3433_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3433_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(5), ack => RPIPE_Block0_start_1320_inst_req_1); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1320_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1323_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1320_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1320_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1323_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1323_Sample/rr
      -- 
    ca_3434_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1320_inst_ack_1, ack => convTransposeA_CP_3352_elements(6)); -- 
    rr_3442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(6), ack => RPIPE_Block0_start_1323_inst_req_0); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1323_Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1323_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1323_Update/cr
      -- CP-element group 7: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1323_update_start_
      -- CP-element group 7: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1323_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1323_Sample/ra
      -- 
    ra_3443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1323_inst_ack_0, ack => convTransposeA_CP_3352_elements(7)); -- 
    cr_3447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(7), ack => RPIPE_Block0_start_1323_inst_req_1); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1326_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1323_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1326_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1323_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1323_Update/ca
      -- CP-element group 8: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1326_Sample/rr
      -- 
    ca_3448_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1323_inst_ack_1, ack => convTransposeA_CP_3352_elements(8)); -- 
    rr_3456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(8), ack => RPIPE_Block0_start_1326_inst_req_0); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1326_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1326_Update/cr
      -- CP-element group 9: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1326_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1326_update_start_
      -- CP-element group 9: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1326_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1326_Sample/$exit
      -- 
    ra_3457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1326_inst_ack_0, ack => convTransposeA_CP_3352_elements(9)); -- 
    cr_3461_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3461_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(9), ack => RPIPE_Block0_start_1326_inst_req_1); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1326_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1329_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1329_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1329_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1326_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1326_Update/$exit
      -- 
    ca_3462_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1326_inst_ack_1, ack => convTransposeA_CP_3352_elements(10)); -- 
    rr_3470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(10), ack => RPIPE_Block0_start_1329_inst_req_0); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1329_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1329_Sample/ra
      -- CP-element group 11: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1329_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1329_update_start_
      -- CP-element group 11: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1329_Update/cr
      -- CP-element group 11: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1329_Update/$entry
      -- 
    ra_3471_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1329_inst_ack_0, ack => convTransposeA_CP_3352_elements(11)); -- 
    cr_3475_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3475_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(11), ack => RPIPE_Block0_start_1329_inst_req_1); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1329_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1329_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1329_Update/ca
      -- CP-element group 12: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1332_sample_start_
      -- CP-element group 12: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1332_Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1332_Sample/rr
      -- 
    ca_3476_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1329_inst_ack_1, ack => convTransposeA_CP_3352_elements(12)); -- 
    rr_3484_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3484_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(12), ack => RPIPE_Block0_start_1332_inst_req_0); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1332_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1332_update_start_
      -- CP-element group 13: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1332_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1332_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1332_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1332_Update/cr
      -- 
    ra_3485_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1332_inst_ack_0, ack => convTransposeA_CP_3352_elements(13)); -- 
    cr_3489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(13), ack => RPIPE_Block0_start_1332_inst_req_1); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1332_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1332_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1332_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1335_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1335_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1335_Sample/rr
      -- 
    ca_3490_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1332_inst_ack_1, ack => convTransposeA_CP_3352_elements(14)); -- 
    rr_3498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(14), ack => RPIPE_Block0_start_1335_inst_req_0); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1335_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1335_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1335_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1335_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1335_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1335_Update/cr
      -- 
    ra_3499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1335_inst_ack_0, ack => convTransposeA_CP_3352_elements(15)); -- 
    cr_3503_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3503_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(15), ack => RPIPE_Block0_start_1335_inst_req_1); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1335_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1335_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1335_Update/ca
      -- CP-element group 16: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1338_sample_start_
      -- CP-element group 16: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1338_Sample/$entry
      -- CP-element group 16: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1338_Sample/rr
      -- 
    ca_3504_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1335_inst_ack_1, ack => convTransposeA_CP_3352_elements(16)); -- 
    rr_3512_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3512_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(16), ack => RPIPE_Block0_start_1338_inst_req_0); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1338_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1338_update_start_
      -- CP-element group 17: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1338_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1338_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1338_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1338_Update/cr
      -- 
    ra_3513_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1338_inst_ack_0, ack => convTransposeA_CP_3352_elements(17)); -- 
    cr_3517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(17), ack => RPIPE_Block0_start_1338_inst_req_1); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1338_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1338_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1338_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1341_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1341_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1341_Sample/rr
      -- 
    ca_3518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1338_inst_ack_1, ack => convTransposeA_CP_3352_elements(18)); -- 
    rr_3526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(18), ack => RPIPE_Block0_start_1341_inst_req_0); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1341_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1341_update_start_
      -- CP-element group 19: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1341_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1341_Sample/ra
      -- CP-element group 19: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1341_Update/$entry
      -- CP-element group 19: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1341_Update/cr
      -- 
    ra_3527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1341_inst_ack_0, ack => convTransposeA_CP_3352_elements(19)); -- 
    cr_3531_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3531_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(19), ack => RPIPE_Block0_start_1341_inst_req_1); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1341_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1341_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1341_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1344_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1344_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1344_Sample/rr
      -- 
    ca_3532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1341_inst_ack_1, ack => convTransposeA_CP_3352_elements(20)); -- 
    rr_3540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(20), ack => RPIPE_Block0_start_1344_inst_req_0); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1344_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1344_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1344_update_start_
      -- CP-element group 21: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1344_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1344_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1344_Update/cr
      -- 
    ra_3541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1344_inst_ack_0, ack => convTransposeA_CP_3352_elements(21)); -- 
    cr_3545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(21), ack => RPIPE_Block0_start_1344_inst_req_1); -- 
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (6) 
      -- CP-element group 22: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1344_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1344_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1344_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1347_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1347_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1347_Sample/rr
      -- 
    ca_3546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1344_inst_ack_1, ack => convTransposeA_CP_3352_elements(22)); -- 
    rr_3554_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3554_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(22), ack => RPIPE_Block0_start_1347_inst_req_0); -- 
    -- CP-element group 23:  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (6) 
      -- CP-element group 23: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1347_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1347_update_start_
      -- CP-element group 23: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1347_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1347_Sample/ra
      -- CP-element group 23: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1347_Update/$entry
      -- CP-element group 23: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1347_Update/cr
      -- 
    ra_3555_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1347_inst_ack_0, ack => convTransposeA_CP_3352_elements(23)); -- 
    cr_3559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(23), ack => RPIPE_Block0_start_1347_inst_req_1); -- 
    -- CP-element group 24:  fork  transition  place  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24: 	26 
    -- CP-element group 24: 	27 
    -- CP-element group 24: 	28 
    -- CP-element group 24: 	29 
    -- CP-element group 24: 	30 
    -- CP-element group 24:  members (25) 
      -- CP-element group 24: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/$exit
      -- CP-element group 24: 	 branch_block_stmt_1312/assign_stmt_1353_to_assign_stmt_1395__entry__
      -- CP-element group 24: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348__exit__
      -- CP-element group 24: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1347_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1347_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_1312/assign_stmt_1315_to_assign_stmt_1348/RPIPE_Block0_start_1347_Update/ca
      -- CP-element group 24: 	 branch_block_stmt_1312/assign_stmt_1353_to_assign_stmt_1395/$entry
      -- CP-element group 24: 	 branch_block_stmt_1312/assign_stmt_1353_to_assign_stmt_1395/type_cast_1352_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1312/assign_stmt_1353_to_assign_stmt_1395/type_cast_1352_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1312/assign_stmt_1353_to_assign_stmt_1395/type_cast_1352_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_1312/assign_stmt_1353_to_assign_stmt_1395/type_cast_1352_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_1312/assign_stmt_1353_to_assign_stmt_1395/type_cast_1352_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1312/assign_stmt_1353_to_assign_stmt_1395/type_cast_1352_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_1312/assign_stmt_1353_to_assign_stmt_1395/type_cast_1356_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1312/assign_stmt_1353_to_assign_stmt_1395/type_cast_1356_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1312/assign_stmt_1353_to_assign_stmt_1395/type_cast_1356_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_1312/assign_stmt_1353_to_assign_stmt_1395/type_cast_1356_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_1312/assign_stmt_1353_to_assign_stmt_1395/type_cast_1356_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1312/assign_stmt_1353_to_assign_stmt_1395/type_cast_1356_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_1312/assign_stmt_1353_to_assign_stmt_1395/type_cast_1366_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1312/assign_stmt_1353_to_assign_stmt_1395/type_cast_1366_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1312/assign_stmt_1353_to_assign_stmt_1395/type_cast_1366_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_1312/assign_stmt_1353_to_assign_stmt_1395/type_cast_1366_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_1312/assign_stmt_1353_to_assign_stmt_1395/type_cast_1366_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1312/assign_stmt_1353_to_assign_stmt_1395/type_cast_1366_Update/cr
      -- 
    ca_3560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1347_inst_ack_1, ack => convTransposeA_CP_3352_elements(24)); -- 
    rr_3571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(24), ack => type_cast_1352_inst_req_0); -- 
    cr_3576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(24), ack => type_cast_1352_inst_req_1); -- 
    rr_3585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(24), ack => type_cast_1356_inst_req_0); -- 
    cr_3590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(24), ack => type_cast_1356_inst_req_1); -- 
    rr_3599_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3599_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(24), ack => type_cast_1366_inst_req_0); -- 
    cr_3604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(24), ack => type_cast_1366_inst_req_1); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_1312/assign_stmt_1353_to_assign_stmt_1395/type_cast_1352_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_1312/assign_stmt_1353_to_assign_stmt_1395/type_cast_1352_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_1312/assign_stmt_1353_to_assign_stmt_1395/type_cast_1352_Sample/ra
      -- 
    ra_3572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1352_inst_ack_0, ack => convTransposeA_CP_3352_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	31 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1312/assign_stmt_1353_to_assign_stmt_1395/type_cast_1352_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_1312/assign_stmt_1353_to_assign_stmt_1395/type_cast_1352_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_1312/assign_stmt_1353_to_assign_stmt_1395/type_cast_1352_Update/ca
      -- 
    ca_3577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1352_inst_ack_1, ack => convTransposeA_CP_3352_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	24 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1312/assign_stmt_1353_to_assign_stmt_1395/type_cast_1356_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_1312/assign_stmt_1353_to_assign_stmt_1395/type_cast_1356_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_1312/assign_stmt_1353_to_assign_stmt_1395/type_cast_1356_Sample/ra
      -- 
    ra_3586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1356_inst_ack_0, ack => convTransposeA_CP_3352_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	24 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	31 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1312/assign_stmt_1353_to_assign_stmt_1395/type_cast_1356_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_1312/assign_stmt_1353_to_assign_stmt_1395/type_cast_1356_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_1312/assign_stmt_1353_to_assign_stmt_1395/type_cast_1356_Update/ca
      -- 
    ca_3591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1356_inst_ack_1, ack => convTransposeA_CP_3352_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	24 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_1312/assign_stmt_1353_to_assign_stmt_1395/type_cast_1366_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_1312/assign_stmt_1353_to_assign_stmt_1395/type_cast_1366_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_1312/assign_stmt_1353_to_assign_stmt_1395/type_cast_1366_Sample/ra
      -- 
    ra_3600_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1366_inst_ack_0, ack => convTransposeA_CP_3352_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	24 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1312/assign_stmt_1353_to_assign_stmt_1395/type_cast_1366_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_1312/assign_stmt_1353_to_assign_stmt_1395/type_cast_1366_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_1312/assign_stmt_1353_to_assign_stmt_1395/type_cast_1366_Update/ca
      -- 
    ca_3605_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1366_inst_ack_1, ack => convTransposeA_CP_3352_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  place  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	26 
    -- CP-element group 31: 	28 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	68 
    -- CP-element group 31: 	69 
    -- CP-element group 31:  members (8) 
      -- CP-element group 31: 	 branch_block_stmt_1312/entry_whilex_xbodyx_xouter
      -- CP-element group 31: 	 branch_block_stmt_1312/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1398/phi_stmt_1398_sources/$entry
      -- CP-element group 31: 	 branch_block_stmt_1312/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1398/$entry
      -- CP-element group 31: 	 branch_block_stmt_1312/assign_stmt_1353_to_assign_stmt_1395__exit__
      -- CP-element group 31: 	 branch_block_stmt_1312/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1405/$entry
      -- CP-element group 31: 	 branch_block_stmt_1312/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1405/phi_stmt_1405_sources/$entry
      -- CP-element group 31: 	 branch_block_stmt_1312/assign_stmt_1353_to_assign_stmt_1395/$exit
      -- CP-element group 31: 	 branch_block_stmt_1312/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- 
    convTransposeA_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3352_elements(26) & convTransposeA_CP_3352_elements(28) & convTransposeA_CP_3352_elements(30);
      gj_convTransposeA_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3352_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	87 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1493_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1493_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1493_Sample/ra
      -- 
    ra_3620_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1493_inst_ack_0, ack => convTransposeA_CP_3352_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	87 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1493_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1493_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1493_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1507_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1507_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1507_Sample/rr
      -- 
    ca_3625_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1493_inst_ack_1, ack => convTransposeA_CP_3352_elements(33)); -- 
    rr_3633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(33), ack => type_cast_1507_inst_req_0); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1507_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1507_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1507_Sample/ra
      -- 
    ra_3634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1507_inst_ack_0, ack => convTransposeA_CP_3352_elements(34)); -- 
    -- CP-element group 35:  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	87 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (16) 
      -- CP-element group 35: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1507_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1507_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1507_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1513_index_resized_1
      -- CP-element group 35: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1513_index_scaled_1
      -- CP-element group 35: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1513_index_computed_1
      -- CP-element group 35: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1513_index_resize_1/$entry
      -- CP-element group 35: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1513_index_resize_1/$exit
      -- CP-element group 35: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1513_index_resize_1/index_resize_req
      -- CP-element group 35: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1513_index_resize_1/index_resize_ack
      -- CP-element group 35: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1513_index_scale_1/$entry
      -- CP-element group 35: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1513_index_scale_1/$exit
      -- CP-element group 35: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1513_index_scale_1/scale_rename_req
      -- CP-element group 35: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1513_index_scale_1/scale_rename_ack
      -- CP-element group 35: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1513_final_index_sum_regn_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1513_final_index_sum_regn_Sample/req
      -- 
    ca_3639_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1507_inst_ack_1, ack => convTransposeA_CP_3352_elements(35)); -- 
    req_3664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(35), ack => array_obj_ref_1513_index_offset_req_0); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	55 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1513_final_index_sum_regn_sample_complete
      -- CP-element group 36: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1513_final_index_sum_regn_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1513_final_index_sum_regn_Sample/ack
      -- 
    ack_3665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1513_index_offset_ack_0, ack => convTransposeA_CP_3352_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	87 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (11) 
      -- CP-element group 37: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/addr_of_1514_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1513_root_address_calculated
      -- CP-element group 37: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1513_offset_calculated
      -- CP-element group 37: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1513_final_index_sum_regn_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1513_final_index_sum_regn_Update/ack
      -- CP-element group 37: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1513_base_plus_offset/$entry
      -- CP-element group 37: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1513_base_plus_offset/$exit
      -- CP-element group 37: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1513_base_plus_offset/sum_rename_req
      -- CP-element group 37: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1513_base_plus_offset/sum_rename_ack
      -- CP-element group 37: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/addr_of_1514_request/$entry
      -- CP-element group 37: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/addr_of_1514_request/req
      -- 
    ack_3670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1513_index_offset_ack_1, ack => convTransposeA_CP_3352_elements(37)); -- 
    req_3679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(37), ack => addr_of_1514_final_reg_req_0); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/addr_of_1514_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/addr_of_1514_request/$exit
      -- CP-element group 38: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/addr_of_1514_request/ack
      -- 
    ack_3680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1514_final_reg_ack_0, ack => convTransposeA_CP_3352_elements(38)); -- 
    -- CP-element group 39:  join  fork  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	87 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (24) 
      -- CP-element group 39: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/addr_of_1514_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/addr_of_1514_complete/$exit
      -- CP-element group 39: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/addr_of_1514_complete/ack
      -- CP-element group 39: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1518_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1518_base_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1518_word_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1518_root_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1518_base_address_resized
      -- CP-element group 39: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1518_base_addr_resize/$entry
      -- CP-element group 39: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1518_base_addr_resize/$exit
      -- CP-element group 39: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1518_base_addr_resize/base_resize_req
      -- CP-element group 39: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1518_base_addr_resize/base_resize_ack
      -- CP-element group 39: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1518_base_plus_offset/$entry
      -- CP-element group 39: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1518_base_plus_offset/$exit
      -- CP-element group 39: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1518_base_plus_offset/sum_rename_req
      -- CP-element group 39: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1518_base_plus_offset/sum_rename_ack
      -- CP-element group 39: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1518_word_addrgen/$entry
      -- CP-element group 39: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1518_word_addrgen/$exit
      -- CP-element group 39: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1518_word_addrgen/root_register_req
      -- CP-element group 39: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1518_word_addrgen/root_register_ack
      -- CP-element group 39: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1518_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1518_Sample/word_access_start/$entry
      -- CP-element group 39: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1518_Sample/word_access_start/word_0/$entry
      -- CP-element group 39: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1518_Sample/word_access_start/word_0/rr
      -- 
    ack_3685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1514_final_reg_ack_1, ack => convTransposeA_CP_3352_elements(39)); -- 
    rr_3718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(39), ack => ptr_deref_1518_load_0_req_0); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (5) 
      -- CP-element group 40: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1518_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1518_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1518_Sample/word_access_start/$exit
      -- CP-element group 40: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1518_Sample/word_access_start/word_0/$exit
      -- CP-element group 40: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1518_Sample/word_access_start/word_0/ra
      -- 
    ra_3719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1518_load_0_ack_0, ack => convTransposeA_CP_3352_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	87 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	50 
    -- CP-element group 41:  members (9) 
      -- CP-element group 41: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1518_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1518_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1518_Update/word_access_complete/$exit
      -- CP-element group 41: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1518_Update/word_access_complete/word_0/$exit
      -- CP-element group 41: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1518_Update/word_access_complete/word_0/ca
      -- CP-element group 41: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1518_Update/ptr_deref_1518_Merge/$entry
      -- CP-element group 41: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1518_Update/ptr_deref_1518_Merge/$exit
      -- CP-element group 41: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1518_Update/ptr_deref_1518_Merge/merge_req
      -- CP-element group 41: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1518_Update/ptr_deref_1518_Merge/merge_ack
      -- 
    ca_3730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1518_load_0_ack_1, ack => convTransposeA_CP_3352_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	87 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1523_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1523_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1523_Sample/ra
      -- 
    ra_3744_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1523_inst_ack_0, ack => convTransposeA_CP_3352_elements(42)); -- 
    -- CP-element group 43:  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	87 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (6) 
      -- CP-element group 43: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1523_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1523_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1523_Update/ca
      -- CP-element group 43: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1537_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1537_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1537_Sample/rr
      -- 
    ca_3749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1523_inst_ack_1, ack => convTransposeA_CP_3352_elements(43)); -- 
    rr_3757_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3757_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(43), ack => type_cast_1537_inst_req_0); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1537_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1537_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1537_Sample/ra
      -- 
    ra_3758_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1537_inst_ack_0, ack => convTransposeA_CP_3352_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	87 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (16) 
      -- CP-element group 45: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1537_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1537_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1537_Update/ca
      -- CP-element group 45: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1543_index_resized_1
      -- CP-element group 45: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1543_index_scaled_1
      -- CP-element group 45: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1543_index_computed_1
      -- CP-element group 45: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1543_index_resize_1/$entry
      -- CP-element group 45: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1543_index_resize_1/$exit
      -- CP-element group 45: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1543_index_resize_1/index_resize_req
      -- CP-element group 45: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1543_index_resize_1/index_resize_ack
      -- CP-element group 45: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1543_index_scale_1/$entry
      -- CP-element group 45: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1543_index_scale_1/$exit
      -- CP-element group 45: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1543_index_scale_1/scale_rename_req
      -- CP-element group 45: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1543_index_scale_1/scale_rename_ack
      -- CP-element group 45: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1543_final_index_sum_regn_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1543_final_index_sum_regn_Sample/req
      -- 
    ca_3763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1537_inst_ack_1, ack => convTransposeA_CP_3352_elements(45)); -- 
    req_3788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(45), ack => array_obj_ref_1543_index_offset_req_0); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	55 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1543_final_index_sum_regn_sample_complete
      -- CP-element group 46: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1543_final_index_sum_regn_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1543_final_index_sum_regn_Sample/ack
      -- 
    ack_3789_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1543_index_offset_ack_0, ack => convTransposeA_CP_3352_elements(46)); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	87 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (11) 
      -- CP-element group 47: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/addr_of_1544_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1543_root_address_calculated
      -- CP-element group 47: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1543_offset_calculated
      -- CP-element group 47: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1543_final_index_sum_regn_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1543_final_index_sum_regn_Update/ack
      -- CP-element group 47: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1543_base_plus_offset/$entry
      -- CP-element group 47: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1543_base_plus_offset/$exit
      -- CP-element group 47: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1543_base_plus_offset/sum_rename_req
      -- CP-element group 47: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1543_base_plus_offset/sum_rename_ack
      -- CP-element group 47: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/addr_of_1544_request/$entry
      -- CP-element group 47: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/addr_of_1544_request/req
      -- 
    ack_3794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1543_index_offset_ack_1, ack => convTransposeA_CP_3352_elements(47)); -- 
    req_3803_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3803_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(47), ack => addr_of_1544_final_reg_req_0); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/addr_of_1544_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/addr_of_1544_request/$exit
      -- CP-element group 48: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/addr_of_1544_request/ack
      -- 
    ack_3804_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1544_final_reg_ack_0, ack => convTransposeA_CP_3352_elements(48)); -- 
    -- CP-element group 49:  fork  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	87 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (19) 
      -- CP-element group 49: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/addr_of_1544_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/addr_of_1544_complete/$exit
      -- CP-element group 49: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/addr_of_1544_complete/ack
      -- CP-element group 49: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1547_base_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1547_word_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1547_root_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1547_base_address_resized
      -- CP-element group 49: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1547_base_addr_resize/$entry
      -- CP-element group 49: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1547_base_addr_resize/$exit
      -- CP-element group 49: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1547_base_addr_resize/base_resize_req
      -- CP-element group 49: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1547_base_addr_resize/base_resize_ack
      -- CP-element group 49: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1547_base_plus_offset/$entry
      -- CP-element group 49: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1547_base_plus_offset/$exit
      -- CP-element group 49: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1547_base_plus_offset/sum_rename_req
      -- CP-element group 49: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1547_base_plus_offset/sum_rename_ack
      -- CP-element group 49: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1547_word_addrgen/$entry
      -- CP-element group 49: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1547_word_addrgen/$exit
      -- CP-element group 49: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1547_word_addrgen/root_register_req
      -- CP-element group 49: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1547_word_addrgen/root_register_ack
      -- 
    ack_3809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1544_final_reg_ack_1, ack => convTransposeA_CP_3352_elements(49)); -- 
    -- CP-element group 50:  join  transition  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	41 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1547_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1547_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1547_Sample/ptr_deref_1547_Split/$entry
      -- CP-element group 50: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1547_Sample/ptr_deref_1547_Split/$exit
      -- CP-element group 50: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1547_Sample/ptr_deref_1547_Split/split_req
      -- CP-element group 50: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1547_Sample/ptr_deref_1547_Split/split_ack
      -- CP-element group 50: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1547_Sample/word_access_start/$entry
      -- CP-element group 50: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1547_Sample/word_access_start/word_0/$entry
      -- CP-element group 50: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1547_Sample/word_access_start/word_0/rr
      -- 
    rr_3847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(50), ack => ptr_deref_1547_store_0_req_0); -- 
    convTransposeA_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3352_elements(41) & convTransposeA_CP_3352_elements(49);
      gj_convTransposeA_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3352_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (5) 
      -- CP-element group 51: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1547_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1547_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1547_Sample/word_access_start/$exit
      -- CP-element group 51: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1547_Sample/word_access_start/word_0/$exit
      -- CP-element group 51: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1547_Sample/word_access_start/word_0/ra
      -- 
    ra_3848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1547_store_0_ack_0, ack => convTransposeA_CP_3352_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	87 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	55 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1547_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1547_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1547_Update/word_access_complete/$exit
      -- CP-element group 52: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1547_Update/word_access_complete/word_0/$exit
      -- CP-element group 52: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1547_Update/word_access_complete/word_0/ca
      -- 
    ca_3859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1547_store_0_ack_1, ack => convTransposeA_CP_3352_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	87 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1553_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1553_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1553_Sample/ra
      -- 
    ra_3868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1553_inst_ack_0, ack => convTransposeA_CP_3352_elements(53)); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	87 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1553_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1553_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1553_Update/ca
      -- 
    ca_3873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1553_inst_ack_1, ack => convTransposeA_CP_3352_elements(54)); -- 
    -- CP-element group 55:  branch  join  transition  place  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	46 
    -- CP-element group 55: 	52 
    -- CP-element group 55: 	54 
    -- CP-element group 55: 	36 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (10) 
      -- CP-element group 55: 	 branch_block_stmt_1312/if_stmt_1568__entry__
      -- CP-element group 55: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567__exit__
      -- CP-element group 55: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/$exit
      -- CP-element group 55: 	 branch_block_stmt_1312/if_stmt_1568_dead_link/$entry
      -- CP-element group 55: 	 branch_block_stmt_1312/if_stmt_1568_eval_test/$entry
      -- CP-element group 55: 	 branch_block_stmt_1312/if_stmt_1568_eval_test/$exit
      -- CP-element group 55: 	 branch_block_stmt_1312/if_stmt_1568_eval_test/branch_req
      -- CP-element group 55: 	 branch_block_stmt_1312/R_cmp_1569_place
      -- CP-element group 55: 	 branch_block_stmt_1312/if_stmt_1568_if_link/$entry
      -- CP-element group 55: 	 branch_block_stmt_1312/if_stmt_1568_else_link/$entry
      -- 
    branch_req_3881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(55), ack => if_stmt_1568_branch_req_0); -- 
    convTransposeA_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3352_elements(46) & convTransposeA_CP_3352_elements(52) & convTransposeA_CP_3352_elements(54) & convTransposeA_CP_3352_elements(36);
      gj_convTransposeA_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3352_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	82 
    -- CP-element group 56: 	83 
    -- CP-element group 56:  members (24) 
      -- CP-element group 56: 	 branch_block_stmt_1312/ifx_xthen_whilex_xbody
      -- CP-element group 56: 	 branch_block_stmt_1312/assign_stmt_1580__entry__
      -- CP-element group 56: 	 branch_block_stmt_1312/merge_stmt_1574__exit__
      -- CP-element group 56: 	 branch_block_stmt_1312/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 56: 	 branch_block_stmt_1312/assign_stmt_1580__exit__
      -- CP-element group 56: 	 branch_block_stmt_1312/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1465/phi_stmt_1465_sources/type_cast_1471/$entry
      -- CP-element group 56: 	 branch_block_stmt_1312/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 56: 	 branch_block_stmt_1312/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1465/$entry
      -- CP-element group 56: 	 branch_block_stmt_1312/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1465/phi_stmt_1465_sources/type_cast_1471/SplitProtocol/Sample/rr
      -- CP-element group 56: 	 branch_block_stmt_1312/merge_stmt_1574_PhiAck/$exit
      -- CP-element group 56: 	 branch_block_stmt_1312/merge_stmt_1574_PhiAck/$entry
      -- CP-element group 56: 	 branch_block_stmt_1312/merge_stmt_1574_PhiReqMerge
      -- CP-element group 56: 	 branch_block_stmt_1312/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1465/phi_stmt_1465_sources/type_cast_1471/SplitProtocol/Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_1312/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1465/phi_stmt_1465_sources/type_cast_1471/SplitProtocol/$entry
      -- CP-element group 56: 	 branch_block_stmt_1312/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 56: 	 branch_block_stmt_1312/merge_stmt_1574_PhiAck/dummy
      -- CP-element group 56: 	 branch_block_stmt_1312/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1465/phi_stmt_1465_sources/$entry
      -- CP-element group 56: 	 branch_block_stmt_1312/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1465/phi_stmt_1465_sources/type_cast_1471/SplitProtocol/Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_1312/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1465/phi_stmt_1465_sources/type_cast_1471/SplitProtocol/Update/cr
      -- CP-element group 56: 	 branch_block_stmt_1312/if_stmt_1568_if_link/$exit
      -- CP-element group 56: 	 branch_block_stmt_1312/if_stmt_1568_if_link/if_choice_transition
      -- CP-element group 56: 	 branch_block_stmt_1312/whilex_xbody_ifx_xthen
      -- CP-element group 56: 	 branch_block_stmt_1312/assign_stmt_1580/$entry
      -- CP-element group 56: 	 branch_block_stmt_1312/assign_stmt_1580/$exit
      -- 
    if_choice_transition_3886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1568_branch_ack_1, ack => convTransposeA_CP_3352_elements(56)); -- 
    rr_4069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(56), ack => type_cast_1471_inst_req_0); -- 
    cr_4074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(56), ack => type_cast_1471_inst_req_1); -- 
    -- CP-element group 57:  fork  transition  place  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57: 	59 
    -- CP-element group 57: 	61 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (24) 
      -- CP-element group 57: 	 branch_block_stmt_1312/merge_stmt_1582__exit__
      -- CP-element group 57: 	 branch_block_stmt_1312/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 57: 	 branch_block_stmt_1312/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 57: 	 branch_block_stmt_1312/assign_stmt_1588_to_assign_stmt_1624/type_cast_1601_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_1312/merge_stmt_1582_PhiReqMerge
      -- CP-element group 57: 	 branch_block_stmt_1312/assign_stmt_1588_to_assign_stmt_1624/type_cast_1601_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_1312/merge_stmt_1582_PhiAck/$entry
      -- CP-element group 57: 	 branch_block_stmt_1312/assign_stmt_1588_to_assign_stmt_1624/type_cast_1618_update_start_
      -- CP-element group 57: 	 branch_block_stmt_1312/assign_stmt_1588_to_assign_stmt_1624__entry__
      -- CP-element group 57: 	 branch_block_stmt_1312/assign_stmt_1588_to_assign_stmt_1624/type_cast_1601_update_start_
      -- CP-element group 57: 	 branch_block_stmt_1312/merge_stmt_1582_PhiAck/$exit
      -- CP-element group 57: 	 branch_block_stmt_1312/merge_stmt_1582_PhiAck/dummy
      -- CP-element group 57: 	 branch_block_stmt_1312/assign_stmt_1588_to_assign_stmt_1624/type_cast_1618_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_1312/assign_stmt_1588_to_assign_stmt_1624/type_cast_1618_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_1312/assign_stmt_1588_to_assign_stmt_1624/type_cast_1592_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_1312/assign_stmt_1588_to_assign_stmt_1624/type_cast_1592_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_1312/if_stmt_1568_else_link/$exit
      -- CP-element group 57: 	 branch_block_stmt_1312/if_stmt_1568_else_link/else_choice_transition
      -- CP-element group 57: 	 branch_block_stmt_1312/whilex_xbody_ifx_xelse
      -- CP-element group 57: 	 branch_block_stmt_1312/assign_stmt_1588_to_assign_stmt_1624/$entry
      -- CP-element group 57: 	 branch_block_stmt_1312/assign_stmt_1588_to_assign_stmt_1624/type_cast_1592_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_1312/assign_stmt_1588_to_assign_stmt_1624/type_cast_1592_update_start_
      -- CP-element group 57: 	 branch_block_stmt_1312/assign_stmt_1588_to_assign_stmt_1624/type_cast_1592_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_1312/assign_stmt_1588_to_assign_stmt_1624/type_cast_1592_Sample/rr
      -- 
    else_choice_transition_3890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1568_branch_ack_0, ack => convTransposeA_CP_3352_elements(57)); -- 
    cr_3925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(57), ack => type_cast_1601_inst_req_1); -- 
    cr_3939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(57), ack => type_cast_1618_inst_req_1); -- 
    cr_3911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(57), ack => type_cast_1592_inst_req_1); -- 
    rr_3906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(57), ack => type_cast_1592_inst_req_0); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_1312/assign_stmt_1588_to_assign_stmt_1624/type_cast_1592_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_1312/assign_stmt_1588_to_assign_stmt_1624/type_cast_1592_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_1312/assign_stmt_1588_to_assign_stmt_1624/type_cast_1592_Sample/ra
      -- 
    ra_3907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1592_inst_ack_0, ack => convTransposeA_CP_3352_elements(58)); -- 
    -- CP-element group 59:  transition  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (6) 
      -- CP-element group 59: 	 branch_block_stmt_1312/assign_stmt_1588_to_assign_stmt_1624/type_cast_1601_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_1312/assign_stmt_1588_to_assign_stmt_1624/type_cast_1601_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_1312/assign_stmt_1588_to_assign_stmt_1624/type_cast_1601_Sample/rr
      -- CP-element group 59: 	 branch_block_stmt_1312/assign_stmt_1588_to_assign_stmt_1624/type_cast_1592_Update/ca
      -- CP-element group 59: 	 branch_block_stmt_1312/assign_stmt_1588_to_assign_stmt_1624/type_cast_1592_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_1312/assign_stmt_1588_to_assign_stmt_1624/type_cast_1592_update_completed_
      -- 
    ca_3912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1592_inst_ack_1, ack => convTransposeA_CP_3352_elements(59)); -- 
    rr_3920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(59), ack => type_cast_1601_inst_req_0); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_1312/assign_stmt_1588_to_assign_stmt_1624/type_cast_1601_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_1312/assign_stmt_1588_to_assign_stmt_1624/type_cast_1601_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_1312/assign_stmt_1588_to_assign_stmt_1624/type_cast_1601_Sample/ra
      -- 
    ra_3921_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1601_inst_ack_0, ack => convTransposeA_CP_3352_elements(60)); -- 
    -- CP-element group 61:  transition  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	57 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_1312/assign_stmt_1588_to_assign_stmt_1624/type_cast_1601_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_1312/assign_stmt_1588_to_assign_stmt_1624/type_cast_1618_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_1312/assign_stmt_1588_to_assign_stmt_1624/type_cast_1601_Update/ca
      -- CP-element group 61: 	 branch_block_stmt_1312/assign_stmt_1588_to_assign_stmt_1624/type_cast_1601_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_1312/assign_stmt_1588_to_assign_stmt_1624/type_cast_1618_Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_1312/assign_stmt_1588_to_assign_stmt_1624/type_cast_1618_Sample/rr
      -- 
    ca_3926_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1601_inst_ack_1, ack => convTransposeA_CP_3352_elements(61)); -- 
    rr_3934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(61), ack => type_cast_1618_inst_req_0); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_1312/assign_stmt_1588_to_assign_stmt_1624/type_cast_1618_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_1312/assign_stmt_1588_to_assign_stmt_1624/type_cast_1618_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_1312/assign_stmt_1588_to_assign_stmt_1624/type_cast_1618_Sample/ra
      -- 
    ra_3935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1618_inst_ack_0, ack => convTransposeA_CP_3352_elements(62)); -- 
    -- CP-element group 63:  branch  transition  place  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (13) 
      -- CP-element group 63: 	 branch_block_stmt_1312/if_stmt_1625_eval_test/$entry
      -- CP-element group 63: 	 branch_block_stmt_1312/assign_stmt_1588_to_assign_stmt_1624/type_cast_1618_Update/ca
      -- CP-element group 63: 	 branch_block_stmt_1312/if_stmt_1625__entry__
      -- CP-element group 63: 	 branch_block_stmt_1312/assign_stmt_1588_to_assign_stmt_1624__exit__
      -- CP-element group 63: 	 branch_block_stmt_1312/if_stmt_1625_eval_test/$exit
      -- CP-element group 63: 	 branch_block_stmt_1312/if_stmt_1625_if_link/$entry
      -- CP-element group 63: 	 branch_block_stmt_1312/if_stmt_1625_eval_test/branch_req
      -- CP-element group 63: 	 branch_block_stmt_1312/assign_stmt_1588_to_assign_stmt_1624/type_cast_1618_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_1312/if_stmt_1625_else_link/$entry
      -- CP-element group 63: 	 branch_block_stmt_1312/assign_stmt_1588_to_assign_stmt_1624/type_cast_1618_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_1312/R_cmp116_1626_place
      -- CP-element group 63: 	 branch_block_stmt_1312/if_stmt_1625_dead_link/$entry
      -- CP-element group 63: 	 branch_block_stmt_1312/assign_stmt_1588_to_assign_stmt_1624/$exit
      -- 
    ca_3940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1618_inst_ack_1, ack => convTransposeA_CP_3352_elements(63)); -- 
    branch_req_3948_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3948_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(63), ack => if_stmt_1625_branch_req_0); -- 
    -- CP-element group 64:  merge  transition  place  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (15) 
      -- CP-element group 64: 	 branch_block_stmt_1312/assign_stmt_1636/$entry
      -- CP-element group 64: 	 branch_block_stmt_1312/ifx_xelse_whilex_xend
      -- CP-element group 64: 	 branch_block_stmt_1312/merge_stmt_1631__exit__
      -- CP-element group 64: 	 branch_block_stmt_1312/assign_stmt_1636__entry__
      -- CP-element group 64: 	 branch_block_stmt_1312/merge_stmt_1631_PhiReqMerge
      -- CP-element group 64: 	 branch_block_stmt_1312/if_stmt_1625_if_link/if_choice_transition
      -- CP-element group 64: 	 branch_block_stmt_1312/if_stmt_1625_if_link/$exit
      -- CP-element group 64: 	 branch_block_stmt_1312/assign_stmt_1636/WPIPE_Block0_done_1633_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_1312/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 64: 	 branch_block_stmt_1312/merge_stmt_1631_PhiAck/$entry
      -- CP-element group 64: 	 branch_block_stmt_1312/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 64: 	 branch_block_stmt_1312/merge_stmt_1631_PhiAck/$exit
      -- CP-element group 64: 	 branch_block_stmt_1312/merge_stmt_1631_PhiAck/dummy
      -- CP-element group 64: 	 branch_block_stmt_1312/assign_stmt_1636/WPIPE_Block0_done_1633_Sample/req
      -- CP-element group 64: 	 branch_block_stmt_1312/assign_stmt_1636/WPIPE_Block0_done_1633_Sample/$entry
      -- 
    if_choice_transition_3953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1625_branch_ack_1, ack => convTransposeA_CP_3352_elements(64)); -- 
    req_3970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(64), ack => WPIPE_Block0_done_1633_inst_req_0); -- 
    -- CP-element group 65:  fork  transition  place  input  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	71 
    -- CP-element group 65: 	72 
    -- CP-element group 65: 	74 
    -- CP-element group 65: 	75 
    -- CP-element group 65:  members (20) 
      -- CP-element group 65: 	 branch_block_stmt_1312/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1405/phi_stmt_1405_sources/type_cast_1411/SplitProtocol/Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1312/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 65: 	 branch_block_stmt_1312/ifx_xelse_whilex_xbodyx_xouter
      -- CP-element group 65: 	 branch_block_stmt_1312/if_stmt_1625_else_link/$exit
      -- CP-element group 65: 	 branch_block_stmt_1312/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1398/$entry
      -- CP-element group 65: 	 branch_block_stmt_1312/if_stmt_1625_else_link/else_choice_transition
      -- CP-element group 65: 	 branch_block_stmt_1312/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1398/phi_stmt_1398_sources/$entry
      -- CP-element group 65: 	 branch_block_stmt_1312/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1405/phi_stmt_1405_sources/type_cast_1411/SplitProtocol/Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1312/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1405/phi_stmt_1405_sources/type_cast_1411/SplitProtocol/Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_1312/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1405/phi_stmt_1405_sources/type_cast_1411/SplitProtocol/Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_1312/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1405/phi_stmt_1405_sources/type_cast_1411/SplitProtocol/$entry
      -- CP-element group 65: 	 branch_block_stmt_1312/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1405/phi_stmt_1405_sources/type_cast_1411/$entry
      -- CP-element group 65: 	 branch_block_stmt_1312/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1405/phi_stmt_1405_sources/$entry
      -- CP-element group 65: 	 branch_block_stmt_1312/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1405/$entry
      -- CP-element group 65: 	 branch_block_stmt_1312/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1398/phi_stmt_1398_sources/type_cast_1404/SplitProtocol/Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1312/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1398/phi_stmt_1398_sources/type_cast_1404/SplitProtocol/Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1312/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1398/phi_stmt_1398_sources/type_cast_1404/SplitProtocol/Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_1312/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1398/phi_stmt_1398_sources/type_cast_1404/SplitProtocol/Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_1312/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1398/phi_stmt_1398_sources/type_cast_1404/SplitProtocol/$entry
      -- CP-element group 65: 	 branch_block_stmt_1312/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1398/phi_stmt_1398_sources/type_cast_1404/$entry
      -- 
    else_choice_transition_3957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1625_branch_ack_0, ack => convTransposeA_CP_3352_elements(65)); -- 
    cr_4042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(65), ack => type_cast_1411_inst_req_1); -- 
    rr_4037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(65), ack => type_cast_1411_inst_req_0); -- 
    cr_4019_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4019_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(65), ack => type_cast_1404_inst_req_1); -- 
    rr_4014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(65), ack => type_cast_1404_inst_req_0); -- 
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_1312/assign_stmt_1636/WPIPE_Block0_done_1633_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_1312/assign_stmt_1636/WPIPE_Block0_done_1633_update_start_
      -- CP-element group 66: 	 branch_block_stmt_1312/assign_stmt_1636/WPIPE_Block0_done_1633_Update/req
      -- CP-element group 66: 	 branch_block_stmt_1312/assign_stmt_1636/WPIPE_Block0_done_1633_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_1312/assign_stmt_1636/WPIPE_Block0_done_1633_Sample/ack
      -- CP-element group 66: 	 branch_block_stmt_1312/assign_stmt_1636/WPIPE_Block0_done_1633_Sample/$exit
      -- 
    ack_3971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1633_inst_ack_0, ack => convTransposeA_CP_3352_elements(66)); -- 
    req_3975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(66), ack => WPIPE_Block0_done_1633_inst_req_1); -- 
    -- CP-element group 67:  transition  place  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (16) 
      -- CP-element group 67: 	 branch_block_stmt_1312/$exit
      -- CP-element group 67: 	 $exit
      -- CP-element group 67: 	 branch_block_stmt_1312/return__
      -- CP-element group 67: 	 branch_block_stmt_1312/assign_stmt_1636__exit__
      -- CP-element group 67: 	 branch_block_stmt_1312/branch_block_stmt_1312__exit__
      -- CP-element group 67: 	 branch_block_stmt_1312/assign_stmt_1636/$exit
      -- CP-element group 67: 	 branch_block_stmt_1312/merge_stmt_1638_PhiReqMerge
      -- CP-element group 67: 	 branch_block_stmt_1312/return___PhiReq/$entry
      -- CP-element group 67: 	 branch_block_stmt_1312/merge_stmt_1638__exit__
      -- CP-element group 67: 	 branch_block_stmt_1312/assign_stmt_1636/WPIPE_Block0_done_1633_Update/ack
      -- CP-element group 67: 	 branch_block_stmt_1312/merge_stmt_1638_PhiAck/dummy
      -- CP-element group 67: 	 branch_block_stmt_1312/merge_stmt_1638_PhiAck/$exit
      -- CP-element group 67: 	 branch_block_stmt_1312/assign_stmt_1636/WPIPE_Block0_done_1633_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_1312/merge_stmt_1638_PhiAck/$entry
      -- CP-element group 67: 	 branch_block_stmt_1312/return___PhiReq/$exit
      -- CP-element group 67: 	 branch_block_stmt_1312/assign_stmt_1636/WPIPE_Block0_done_1633_update_completed_
      -- 
    ack_3976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1633_inst_ack_1, ack => convTransposeA_CP_3352_elements(67)); -- 
    -- CP-element group 68:  transition  output  delay-element  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	31 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (4) 
      -- CP-element group 68: 	 branch_block_stmt_1312/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1398/$exit
      -- CP-element group 68: 	 branch_block_stmt_1312/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1398/phi_stmt_1398_sources/type_cast_1402_konst_delay_trans
      -- CP-element group 68: 	 branch_block_stmt_1312/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1398/phi_stmt_1398_sources/$exit
      -- CP-element group 68: 	 branch_block_stmt_1312/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1398/phi_stmt_1398_req
      -- 
    phi_stmt_1398_req_3987_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1398_req_3987_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(68), ack => phi_stmt_1398_req_0); -- 
    -- Element group convTransposeA_CP_3352_elements(68) is a control-delay.
    cp_element_68_delay: control_delay_element  generic map(name => " 68_delay", delay_value => 1)  port map(req => convTransposeA_CP_3352_elements(31), ack => convTransposeA_CP_3352_elements(68), clk => clk, reset =>reset);
    -- CP-element group 69:  transition  output  delay-element  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	31 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (4) 
      -- CP-element group 69: 	 branch_block_stmt_1312/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1405/phi_stmt_1405_sources/type_cast_1409_konst_delay_trans
      -- CP-element group 69: 	 branch_block_stmt_1312/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1405/phi_stmt_1405_req
      -- CP-element group 69: 	 branch_block_stmt_1312/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1405/phi_stmt_1405_sources/$exit
      -- CP-element group 69: 	 branch_block_stmt_1312/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1405/$exit
      -- 
    phi_stmt_1405_req_3995_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1405_req_3995_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(69), ack => phi_stmt_1405_req_0); -- 
    -- Element group convTransposeA_CP_3352_elements(69) is a control-delay.
    cp_element_69_delay: control_delay_element  generic map(name => " 69_delay", delay_value => 1)  port map(req => convTransposeA_CP_3352_elements(31), ack => convTransposeA_CP_3352_elements(69), clk => clk, reset =>reset);
    -- CP-element group 70:  join  transition  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	78 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_1312/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3352_elements(68) & convTransposeA_CP_3352_elements(69);
      gj_convTransposeA_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3352_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	65 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (2) 
      -- CP-element group 71: 	 branch_block_stmt_1312/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1398/phi_stmt_1398_sources/type_cast_1404/SplitProtocol/Sample/ra
      -- CP-element group 71: 	 branch_block_stmt_1312/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1398/phi_stmt_1398_sources/type_cast_1404/SplitProtocol/Sample/$exit
      -- 
    ra_4015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1404_inst_ack_0, ack => convTransposeA_CP_3352_elements(71)); -- 
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	65 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (2) 
      -- CP-element group 72: 	 branch_block_stmt_1312/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1398/phi_stmt_1398_sources/type_cast_1404/SplitProtocol/Update/ca
      -- CP-element group 72: 	 branch_block_stmt_1312/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1398/phi_stmt_1398_sources/type_cast_1404/SplitProtocol/Update/$exit
      -- 
    ca_4020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1404_inst_ack_1, ack => convTransposeA_CP_3352_elements(72)); -- 
    -- CP-element group 73:  join  transition  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	77 
    -- CP-element group 73:  members (5) 
      -- CP-element group 73: 	 branch_block_stmt_1312/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1398/$exit
      -- CP-element group 73: 	 branch_block_stmt_1312/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1398/phi_stmt_1398_req
      -- CP-element group 73: 	 branch_block_stmt_1312/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1398/phi_stmt_1398_sources/type_cast_1404/SplitProtocol/$exit
      -- CP-element group 73: 	 branch_block_stmt_1312/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1398/phi_stmt_1398_sources/type_cast_1404/$exit
      -- CP-element group 73: 	 branch_block_stmt_1312/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1398/phi_stmt_1398_sources/$exit
      -- 
    phi_stmt_1398_req_4021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1398_req_4021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(73), ack => phi_stmt_1398_req_1); -- 
    convTransposeA_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3352_elements(71) & convTransposeA_CP_3352_elements(72);
      gj_convTransposeA_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3352_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	65 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (2) 
      -- CP-element group 74: 	 branch_block_stmt_1312/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1405/phi_stmt_1405_sources/type_cast_1411/SplitProtocol/Sample/ra
      -- CP-element group 74: 	 branch_block_stmt_1312/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1405/phi_stmt_1405_sources/type_cast_1411/SplitProtocol/Sample/$exit
      -- 
    ra_4038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1411_inst_ack_0, ack => convTransposeA_CP_3352_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	65 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_1312/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1405/phi_stmt_1405_sources/type_cast_1411/SplitProtocol/Update/ca
      -- CP-element group 75: 	 branch_block_stmt_1312/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1405/phi_stmt_1405_sources/type_cast_1411/SplitProtocol/Update/$exit
      -- 
    ca_4043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1411_inst_ack_1, ack => convTransposeA_CP_3352_elements(75)); -- 
    -- CP-element group 76:  join  transition  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (5) 
      -- CP-element group 76: 	 branch_block_stmt_1312/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1405/phi_stmt_1405_req
      -- CP-element group 76: 	 branch_block_stmt_1312/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1405/phi_stmt_1405_sources/type_cast_1411/SplitProtocol/$exit
      -- CP-element group 76: 	 branch_block_stmt_1312/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1405/phi_stmt_1405_sources/type_cast_1411/$exit
      -- CP-element group 76: 	 branch_block_stmt_1312/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1405/phi_stmt_1405_sources/$exit
      -- CP-element group 76: 	 branch_block_stmt_1312/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1405/$exit
      -- 
    phi_stmt_1405_req_4044_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1405_req_4044_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(76), ack => phi_stmt_1405_req_1); -- 
    convTransposeA_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3352_elements(74) & convTransposeA_CP_3352_elements(75);
      gj_convTransposeA_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3352_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  join  transition  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	73 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_1312/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3352_elements(73) & convTransposeA_CP_3352_elements(76);
      gj_convTransposeA_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3352_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  merge  fork  transition  place  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	70 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (2) 
      -- CP-element group 78: 	 branch_block_stmt_1312/merge_stmt_1397_PhiAck/$entry
      -- CP-element group 78: 	 branch_block_stmt_1312/merge_stmt_1397_PhiReqMerge
      -- 
    convTransposeA_CP_3352_elements(78) <= OrReduce(convTransposeA_CP_3352_elements(70) & convTransposeA_CP_3352_elements(77));
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_1312/merge_stmt_1397_PhiAck/phi_stmt_1398_ack
      -- 
    phi_stmt_1398_ack_4049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1398_ack_0, ack => convTransposeA_CP_3352_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_1312/merge_stmt_1397_PhiAck/phi_stmt_1405_ack
      -- 
    phi_stmt_1405_ack_4050_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1405_ack_0, ack => convTransposeA_CP_3352_elements(80)); -- 
    -- CP-element group 81:  join  transition  place  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	85 
    -- CP-element group 81:  members (10) 
      -- CP-element group 81: 	 branch_block_stmt_1312/assign_stmt_1417_to_assign_stmt_1462__exit__
      -- CP-element group 81: 	 branch_block_stmt_1312/merge_stmt_1397__exit__
      -- CP-element group 81: 	 branch_block_stmt_1312/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 81: 	 branch_block_stmt_1312/merge_stmt_1397_PhiAck/$exit
      -- CP-element group 81: 	 branch_block_stmt_1312/assign_stmt_1417_to_assign_stmt_1462__entry__
      -- CP-element group 81: 	 branch_block_stmt_1312/assign_stmt_1417_to_assign_stmt_1462/$entry
      -- CP-element group 81: 	 branch_block_stmt_1312/assign_stmt_1417_to_assign_stmt_1462/$exit
      -- CP-element group 81: 	 branch_block_stmt_1312/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1465/phi_stmt_1465_sources/$entry
      -- CP-element group 81: 	 branch_block_stmt_1312/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1465/$entry
      -- CP-element group 81: 	 branch_block_stmt_1312/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- 
    convTransposeA_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3352_elements(79) & convTransposeA_CP_3352_elements(80);
      gj_convTransposeA_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3352_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	56 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_1312/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1465/phi_stmt_1465_sources/type_cast_1471/SplitProtocol/Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_1312/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1465/phi_stmt_1465_sources/type_cast_1471/SplitProtocol/Sample/ra
      -- 
    ra_4070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1471_inst_ack_0, ack => convTransposeA_CP_3352_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	56 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_1312/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1465/phi_stmt_1465_sources/type_cast_1471/SplitProtocol/Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_1312/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1465/phi_stmt_1465_sources/type_cast_1471/SplitProtocol/Update/ca
      -- 
    ca_4075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1471_inst_ack_1, ack => convTransposeA_CP_3352_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (6) 
      -- CP-element group 84: 	 branch_block_stmt_1312/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1465/$exit
      -- CP-element group 84: 	 branch_block_stmt_1312/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- CP-element group 84: 	 branch_block_stmt_1312/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1465/phi_stmt_1465_sources/type_cast_1471/$exit
      -- CP-element group 84: 	 branch_block_stmt_1312/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1465/phi_stmt_1465_sources/type_cast_1471/SplitProtocol/$exit
      -- CP-element group 84: 	 branch_block_stmt_1312/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1465/phi_stmt_1465_sources/$exit
      -- CP-element group 84: 	 branch_block_stmt_1312/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1465/phi_stmt_1465_req
      -- 
    phi_stmt_1465_req_4076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1465_req_4076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(84), ack => phi_stmt_1465_req_1); -- 
    convTransposeA_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3352_elements(82) & convTransposeA_CP_3352_elements(83);
      gj_convTransposeA_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3352_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  transition  output  delay-element  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	81 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (5) 
      -- CP-element group 85: 	 branch_block_stmt_1312/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1465/phi_stmt_1465_req
      -- CP-element group 85: 	 branch_block_stmt_1312/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1465/phi_stmt_1465_sources/type_cast_1469_konst_delay_trans
      -- CP-element group 85: 	 branch_block_stmt_1312/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1465/phi_stmt_1465_sources/$exit
      -- CP-element group 85: 	 branch_block_stmt_1312/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1465/$exit
      -- CP-element group 85: 	 branch_block_stmt_1312/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- 
    phi_stmt_1465_req_4087_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1465_req_4087_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(85), ack => phi_stmt_1465_req_0); -- 
    -- Element group convTransposeA_CP_3352_elements(85) is a control-delay.
    cp_element_85_delay: control_delay_element  generic map(name => " 85_delay", delay_value => 1)  port map(req => convTransposeA_CP_3352_elements(81), ack => convTransposeA_CP_3352_elements(85), clk => clk, reset =>reset);
    -- CP-element group 86:  merge  transition  place  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_1312/merge_stmt_1464_PhiReqMerge
      -- CP-element group 86: 	 branch_block_stmt_1312/merge_stmt_1464_PhiAck/$entry
      -- 
    convTransposeA_CP_3352_elements(86) <= OrReduce(convTransposeA_CP_3352_elements(84) & convTransposeA_CP_3352_elements(85));
    -- CP-element group 87:  fork  transition  place  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	41 
    -- CP-element group 87: 	42 
    -- CP-element group 87: 	43 
    -- CP-element group 87: 	45 
    -- CP-element group 87: 	47 
    -- CP-element group 87: 	49 
    -- CP-element group 87: 	52 
    -- CP-element group 87: 	53 
    -- CP-element group 87: 	54 
    -- CP-element group 87: 	32 
    -- CP-element group 87: 	33 
    -- CP-element group 87: 	35 
    -- CP-element group 87: 	37 
    -- CP-element group 87: 	39 
    -- CP-element group 87:  members (51) 
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567__entry__
      -- CP-element group 87: 	 branch_block_stmt_1312/merge_stmt_1464__exit__
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/$entry
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1493_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1493_update_start_
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1493_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1493_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_1312/merge_stmt_1464_PhiAck/phi_stmt_1465_ack
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1493_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1493_Update/cr
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1507_update_start_
      -- CP-element group 87: 	 branch_block_stmt_1312/merge_stmt_1464_PhiAck/$exit
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1507_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1507_Update/cr
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/addr_of_1514_update_start_
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1513_final_index_sum_regn_update_start
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1513_final_index_sum_regn_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1513_final_index_sum_regn_Update/req
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/addr_of_1514_complete/$entry
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/addr_of_1514_complete/req
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1518_update_start_
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1518_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1518_Update/word_access_complete/$entry
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1518_Update/word_access_complete/word_0/$entry
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1518_Update/word_access_complete/word_0/cr
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1523_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1523_update_start_
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1523_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1523_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1523_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1523_Update/cr
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1537_update_start_
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1537_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1537_Update/cr
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/addr_of_1544_update_start_
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1543_final_index_sum_regn_update_start
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1543_final_index_sum_regn_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/array_obj_ref_1543_final_index_sum_regn_Update/req
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/addr_of_1544_complete/$entry
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/addr_of_1544_complete/req
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1547_update_start_
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1547_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1547_Update/word_access_complete/$entry
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1547_Update/word_access_complete/word_0/$entry
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/ptr_deref_1547_Update/word_access_complete/word_0/cr
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1553_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1553_update_start_
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1553_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1553_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1553_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_1312/assign_stmt_1478_to_assign_stmt_1567/type_cast_1553_Update/cr
      -- 
    phi_stmt_1465_ack_4092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1465_ack_0, ack => convTransposeA_CP_3352_elements(87)); -- 
    rr_3619_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3619_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(87), ack => type_cast_1493_inst_req_0); -- 
    cr_3624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(87), ack => type_cast_1493_inst_req_1); -- 
    cr_3638_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3638_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(87), ack => type_cast_1507_inst_req_1); -- 
    req_3669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(87), ack => array_obj_ref_1513_index_offset_req_1); -- 
    req_3684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(87), ack => addr_of_1514_final_reg_req_1); -- 
    cr_3729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(87), ack => ptr_deref_1518_load_0_req_1); -- 
    rr_3743_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3743_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(87), ack => type_cast_1523_inst_req_0); -- 
    cr_3748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(87), ack => type_cast_1523_inst_req_1); -- 
    cr_3762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(87), ack => type_cast_1537_inst_req_1); -- 
    req_3793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(87), ack => array_obj_ref_1543_index_offset_req_1); -- 
    req_3808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(87), ack => addr_of_1544_final_reg_req_1); -- 
    cr_3858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(87), ack => ptr_deref_1547_store_0_req_1); -- 
    rr_3867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(87), ack => type_cast_1553_inst_req_0); -- 
    cr_3872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3352_elements(87), ack => type_cast_1553_inst_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_1501_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1531_wire : std_logic_vector(31 downto 0);
    signal R_idxprom85_1542_resized : std_logic_vector(13 downto 0);
    signal R_idxprom85_1542_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_1512_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_1512_scaled : std_logic_vector(13 downto 0);
    signal add32_1483 : std_logic_vector(15 downto 0);
    signal add76_1488 : std_logic_vector(15 downto 0);
    signal add90_1560 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1513_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1513_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1513_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1513_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1513_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1513_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1543_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1543_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1543_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1543_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1543_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1543_root_address : std_logic_vector(13 downto 0);
    signal arrayidx80_1515 : std_logic_vector(31 downto 0);
    signal arrayidx86_1545 : std_logic_vector(31 downto 0);
    signal call11_1333 : std_logic_vector(15 downto 0);
    signal call13_1336 : std_logic_vector(15 downto 0);
    signal call14_1339 : std_logic_vector(15 downto 0);
    signal call15_1342 : std_logic_vector(15 downto 0);
    signal call17_1345 : std_logic_vector(15 downto 0);
    signal call19_1348 : std_logic_vector(15 downto 0);
    signal call1_1318 : std_logic_vector(15 downto 0);
    signal call3_1321 : std_logic_vector(15 downto 0);
    signal call5_1324 : std_logic_vector(15 downto 0);
    signal call7_1327 : std_logic_vector(15 downto 0);
    signal call9_1330 : std_logic_vector(15 downto 0);
    signal call_1315 : std_logic_vector(15 downto 0);
    signal cmp105_1598 : std_logic_vector(0 downto 0);
    signal cmp116_1624 : std_logic_vector(0 downto 0);
    signal cmp_1567 : std_logic_vector(0 downto 0);
    signal conv101_1593 : std_logic_vector(31 downto 0);
    signal conv104_1357 : std_logic_vector(31 downto 0);
    signal conv111_1619 : std_logic_vector(31 downto 0);
    signal conv114_1367 : std_logic_vector(31 downto 0);
    signal conv79_1494 : std_logic_vector(31 downto 0);
    signal conv83_1524 : std_logic_vector(31 downto 0);
    signal conv89_1554 : std_logic_vector(31 downto 0);
    signal conv93_1353 : std_logic_vector(31 downto 0);
    signal div115_1373 : std_logic_vector(31 downto 0);
    signal div_1363 : std_logic_vector(31 downto 0);
    signal idxprom85_1538 : std_logic_vector(63 downto 0);
    signal idxprom_1508 : std_logic_vector(63 downto 0);
    signal inc109_1602 : std_logic_vector(15 downto 0);
    signal inc109x_xinput_dim0x_x2_1607 : std_logic_vector(15 downto 0);
    signal inc_1588 : std_logic_vector(15 downto 0);
    signal indvar_1465 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_1580 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_1405 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_1398 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_1614 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1478 : std_logic_vector(15 downto 0);
    signal ptr_deref_1518_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1518_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1518_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1518_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1518_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1547_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1547_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1547_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1547_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1547_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1547_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr84_1533 : std_logic_vector(31 downto 0);
    signal shr_1503 : std_logic_vector(31 downto 0);
    signal tmp10_1462 : std_logic_vector(15 downto 0);
    signal tmp143_1417 : std_logic_vector(15 downto 0);
    signal tmp144_1422 : std_logic_vector(15 downto 0);
    signal tmp145_1427 : std_logic_vector(15 downto 0);
    signal tmp1_1384 : std_logic_vector(15 downto 0);
    signal tmp2_1432 : std_logic_vector(15 downto 0);
    signal tmp3_1437 : std_logic_vector(15 downto 0);
    signal tmp4_1390 : std_logic_vector(15 downto 0);
    signal tmp5_1395 : std_logic_vector(15 downto 0);
    signal tmp6_1442 : std_logic_vector(15 downto 0);
    signal tmp7_1447 : std_logic_vector(15 downto 0);
    signal tmp81_1519 : std_logic_vector(63 downto 0);
    signal tmp8_1452 : std_logic_vector(15 downto 0);
    signal tmp9_1457 : std_logic_vector(15 downto 0);
    signal tmp_1379 : std_logic_vector(15 downto 0);
    signal type_cast_1361_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1371_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1377_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1388_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1402_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1404_wire : std_logic_vector(15 downto 0);
    signal type_cast_1409_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1411_wire : std_logic_vector(15 downto 0);
    signal type_cast_1469_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1471_wire : std_logic_vector(15 downto 0);
    signal type_cast_1476_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1492_wire : std_logic_vector(31 downto 0);
    signal type_cast_1497_wire : std_logic_vector(31 downto 0);
    signal type_cast_1500_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1506_wire : std_logic_vector(63 downto 0);
    signal type_cast_1522_wire : std_logic_vector(31 downto 0);
    signal type_cast_1527_wire : std_logic_vector(31 downto 0);
    signal type_cast_1530_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1536_wire : std_logic_vector(63 downto 0);
    signal type_cast_1552_wire : std_logic_vector(31 downto 0);
    signal type_cast_1558_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1563_wire : std_logic_vector(31 downto 0);
    signal type_cast_1565_wire : std_logic_vector(31 downto 0);
    signal type_cast_1578_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1586_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1591_wire : std_logic_vector(31 downto 0);
    signal type_cast_1611_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1617_wire : std_logic_vector(31 downto 0);
    signal type_cast_1635_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_1513_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1513_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1513_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1513_resized_base_address <= "00000000000000";
    array_obj_ref_1543_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1543_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1543_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1543_resized_base_address <= "00000000000000";
    ptr_deref_1518_word_offset_0 <= "00000000000000";
    ptr_deref_1547_word_offset_0 <= "00000000000000";
    type_cast_1361_wire_constant <= "00000000000000000000000000000001";
    type_cast_1371_wire_constant <= "00000000000000000000000000000001";
    type_cast_1377_wire_constant <= "1111111111111111";
    type_cast_1388_wire_constant <= "1111111111111111";
    type_cast_1402_wire_constant <= "0000000000000000";
    type_cast_1409_wire_constant <= "0000000000000000";
    type_cast_1469_wire_constant <= "0000000000000000";
    type_cast_1476_wire_constant <= "0000000000000100";
    type_cast_1500_wire_constant <= "00000000000000000000000000000010";
    type_cast_1530_wire_constant <= "00000000000000000000000000000010";
    type_cast_1558_wire_constant <= "00000000000000000000000000000100";
    type_cast_1578_wire_constant <= "0000000000000001";
    type_cast_1586_wire_constant <= "0000000000000001";
    type_cast_1611_wire_constant <= "0000000000000000";
    type_cast_1635_wire_constant <= "0000000000000001";
    phi_stmt_1398: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1402_wire_constant & type_cast_1404_wire;
      req <= phi_stmt_1398_req_0 & phi_stmt_1398_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1398",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1398_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_1398,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1398
    phi_stmt_1405: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1409_wire_constant & type_cast_1411_wire;
      req <= phi_stmt_1405_req_0 & phi_stmt_1405_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1405",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1405_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_1405,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1405
    phi_stmt_1465: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1469_wire_constant & type_cast_1471_wire;
      req <= phi_stmt_1465_req_0 & phi_stmt_1465_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1465",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1465_ack_0,
          idata => idata,
          odata => indvar_1465,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1465
    -- flow-through select operator MUX_1613_inst
    input_dim1x_x2_1614 <= type_cast_1611_wire_constant when (cmp105_1598(0) /=  '0') else inc_1588;
    addr_of_1514_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1514_final_reg_req_0;
      addr_of_1514_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1514_final_reg_req_1;
      addr_of_1514_final_reg_ack_1<= rack(0);
      addr_of_1514_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1514_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1513_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx80_1515,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1544_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1544_final_reg_req_0;
      addr_of_1544_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1544_final_reg_req_1;
      addr_of_1544_final_reg_ack_1<= rack(0);
      addr_of_1544_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1544_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1543_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx86_1545,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1352_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1352_inst_req_0;
      type_cast_1352_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1352_inst_req_1;
      type_cast_1352_inst_ack_1<= rack(0);
      type_cast_1352_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1352_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_1321,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv93_1353,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1356_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1356_inst_req_0;
      type_cast_1356_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1356_inst_req_1;
      type_cast_1356_inst_ack_1<= rack(0);
      type_cast_1356_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1356_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1_1318,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv104_1357,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1366_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1366_inst_req_0;
      type_cast_1366_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1366_inst_req_1;
      type_cast_1366_inst_ack_1<= rack(0);
      type_cast_1366_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1366_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1315,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv114_1367,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1404_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1404_inst_req_0;
      type_cast_1404_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1404_inst_req_1;
      type_cast_1404_inst_ack_1<= rack(0);
      type_cast_1404_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1404_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_1614,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1404_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1411_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1411_inst_req_0;
      type_cast_1411_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1411_inst_req_1;
      type_cast_1411_inst_ack_1<= rack(0);
      type_cast_1411_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1411_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc109x_xinput_dim0x_x2_1607,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1411_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1471_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1471_inst_req_0;
      type_cast_1471_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1471_inst_req_1;
      type_cast_1471_inst_ack_1<= rack(0);
      type_cast_1471_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1471_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1580,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1471_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1493_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1493_inst_req_0;
      type_cast_1493_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1493_inst_req_1;
      type_cast_1493_inst_ack_1<= rack(0);
      type_cast_1493_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1493_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1492_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv79_1494,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1497_inst
    process(conv79_1494) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv79_1494(31 downto 0);
      type_cast_1497_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1502_inst
    process(ASHR_i32_i32_1501_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1501_wire(31 downto 0);
      shr_1503 <= tmp_var; -- 
    end process;
    type_cast_1507_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1507_inst_req_0;
      type_cast_1507_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1507_inst_req_1;
      type_cast_1507_inst_ack_1<= rack(0);
      type_cast_1507_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1507_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1506_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_1508,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1523_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1523_inst_req_0;
      type_cast_1523_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1523_inst_req_1;
      type_cast_1523_inst_ack_1<= rack(0);
      type_cast_1523_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1523_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1522_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv83_1524,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1527_inst
    process(conv83_1524) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv83_1524(31 downto 0);
      type_cast_1527_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1532_inst
    process(ASHR_i32_i32_1531_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1531_wire(31 downto 0);
      shr84_1533 <= tmp_var; -- 
    end process;
    type_cast_1537_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1537_inst_req_0;
      type_cast_1537_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1537_inst_req_1;
      type_cast_1537_inst_ack_1<= rack(0);
      type_cast_1537_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1537_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1536_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom85_1538,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1553_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1553_inst_req_0;
      type_cast_1553_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1553_inst_req_1;
      type_cast_1553_inst_ack_1<= rack(0);
      type_cast_1553_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1553_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1552_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv89_1554,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1563_inst
    process(add90_1560) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add90_1560(31 downto 0);
      type_cast_1563_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1565_inst
    process(conv93_1353) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv93_1353(31 downto 0);
      type_cast_1565_wire <= tmp_var; -- 
    end process;
    type_cast_1592_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1592_inst_req_0;
      type_cast_1592_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1592_inst_req_1;
      type_cast_1592_inst_ack_1<= rack(0);
      type_cast_1592_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1592_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1591_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv101_1593,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1601_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1601_inst_req_0;
      type_cast_1601_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1601_inst_req_1;
      type_cast_1601_inst_ack_1<= rack(0);
      type_cast_1601_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1601_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp105_1598,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc109_1602,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1618_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1618_inst_req_0;
      type_cast_1618_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1618_inst_req_1;
      type_cast_1618_inst_ack_1<= rack(0);
      type_cast_1618_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1618_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1617_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv111_1619,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1513_index_1_rename
    process(R_idxprom_1512_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_1512_resized;
      ov(13 downto 0) := iv;
      R_idxprom_1512_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1513_index_1_resize
    process(idxprom_1508) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_1508;
      ov := iv(13 downto 0);
      R_idxprom_1512_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1513_root_address_inst
    process(array_obj_ref_1513_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1513_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1513_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1543_index_1_rename
    process(R_idxprom85_1542_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom85_1542_resized;
      ov(13 downto 0) := iv;
      R_idxprom85_1542_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1543_index_1_resize
    process(idxprom85_1538) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom85_1538;
      ov := iv(13 downto 0);
      R_idxprom85_1542_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1543_root_address_inst
    process(array_obj_ref_1543_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1543_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1543_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1518_addr_0
    process(ptr_deref_1518_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1518_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1518_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1518_base_resize
    process(arrayidx80_1515) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx80_1515;
      ov := iv(13 downto 0);
      ptr_deref_1518_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1518_gather_scatter
    process(ptr_deref_1518_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1518_data_0;
      ov(63 downto 0) := iv;
      tmp81_1519 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1518_root_address_inst
    process(ptr_deref_1518_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1518_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1518_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1547_addr_0
    process(ptr_deref_1547_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1547_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1547_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1547_base_resize
    process(arrayidx86_1545) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx86_1545;
      ov := iv(13 downto 0);
      ptr_deref_1547_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1547_gather_scatter
    process(tmp81_1519) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp81_1519;
      ov(63 downto 0) := iv;
      ptr_deref_1547_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1547_root_address_inst
    process(ptr_deref_1547_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1547_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1547_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1568_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_1567;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1568_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1568_branch_req_0,
          ack0 => if_stmt_1568_branch_ack_0,
          ack1 => if_stmt_1568_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1625_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp116_1624;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1625_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1625_branch_req_0,
          ack0 => if_stmt_1625_branch_ack_0,
          ack1 => if_stmt_1625_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1378_inst
    process(call9_1330) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_1330, type_cast_1377_wire_constant, tmp_var);
      tmp_1379 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1389_inst
    process(call7_1327) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_1327, type_cast_1388_wire_constant, tmp_var);
      tmp4_1390 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1421_inst
    process(input_dim1x_x1x_xph_1398, tmp143_1417) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_1398, tmp143_1417, tmp_var);
      tmp144_1422 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1436_inst
    process(tmp1_1384, tmp2_1432) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp1_1384, tmp2_1432, tmp_var);
      tmp3_1437 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1446_inst
    process(tmp5_1395, tmp6_1442) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp5_1395, tmp6_1442, tmp_var);
      tmp7_1447 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1456_inst
    process(tmp3_1437, tmp8_1452) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp3_1437, tmp8_1452, tmp_var);
      tmp9_1457 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1482_inst
    process(tmp145_1427, input_dim2x_x1_1478) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp145_1427, input_dim2x_x1_1478, tmp_var);
      add32_1483 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1487_inst
    process(tmp10_1462, input_dim2x_x1_1478) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp10_1462, input_dim2x_x1_1478, tmp_var);
      add76_1488 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1579_inst
    process(indvar_1465) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1465, type_cast_1578_wire_constant, tmp_var);
      indvarx_xnext_1580 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1587_inst
    process(input_dim1x_x1x_xph_1398) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_1398, type_cast_1586_wire_constant, tmp_var);
      inc_1588 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1606_inst
    process(inc109_1602, input_dim0x_x2x_xph_1405) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc109_1602, input_dim0x_x2x_xph_1405, tmp_var);
      inc109x_xinput_dim0x_x2_1607 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1559_inst
    process(conv89_1554) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv89_1554, type_cast_1558_wire_constant, tmp_var);
      add90_1560 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1501_inst
    process(type_cast_1497_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1497_wire, type_cast_1500_wire_constant, tmp_var);
      ASHR_i32_i32_1501_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1531_inst
    process(type_cast_1527_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1527_wire, type_cast_1530_wire_constant, tmp_var);
      ASHR_i32_i32_1531_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1597_inst
    process(conv101_1593, div_1363) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv101_1593, div_1363, tmp_var);
      cmp105_1598 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1623_inst
    process(conv111_1619, div115_1373) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv111_1619, div115_1373, tmp_var);
      cmp116_1624 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1362_inst
    process(conv104_1357) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv104_1357, type_cast_1361_wire_constant, tmp_var);
      div_1363 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1372_inst
    process(conv114_1367) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv114_1367, type_cast_1371_wire_constant, tmp_var);
      div115_1373 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1416_inst
    process(call1_1318, input_dim0x_x2x_xph_1405) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call1_1318, input_dim0x_x2x_xph_1405, tmp_var);
      tmp143_1417 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1426_inst
    process(call3_1321, tmp144_1422) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call3_1321, tmp144_1422, tmp_var);
      tmp145_1427 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1431_inst
    process(call13_1336, input_dim1x_x1x_xph_1398) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call13_1336, input_dim1x_x1x_xph_1398, tmp_var);
      tmp2_1432 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1441_inst
    process(call13_1336, input_dim0x_x2x_xph_1405) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call13_1336, input_dim0x_x2x_xph_1405, tmp_var);
      tmp6_1442 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1451_inst
    process(call17_1345, tmp7_1447) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call17_1345, tmp7_1447, tmp_var);
      tmp8_1452 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1461_inst
    process(call19_1348, tmp9_1457) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call19_1348, tmp9_1457, tmp_var);
      tmp10_1462 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1477_inst
    process(indvar_1465) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_1465, type_cast_1476_wire_constant, tmp_var);
      input_dim2x_x1_1478 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1566_inst
    process(type_cast_1563_wire, type_cast_1565_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1563_wire, type_cast_1565_wire, tmp_var);
      cmp_1567 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1383_inst
    process(tmp_1379, call14_1339) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp_1379, call14_1339, tmp_var);
      tmp1_1384 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1394_inst
    process(tmp4_1390, call14_1339) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp4_1390, call14_1339, tmp_var);
      tmp5_1395 <= tmp_var; --
    end process;
    -- shared split operator group (28) : array_obj_ref_1513_index_offset 
    ApIntAdd_group_28: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_1512_scaled;
      array_obj_ref_1513_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1513_index_offset_req_0;
      array_obj_ref_1513_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1513_index_offset_req_1;
      array_obj_ref_1513_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_28_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_28_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : array_obj_ref_1543_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom85_1542_scaled;
      array_obj_ref_1543_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1543_index_offset_req_0;
      array_obj_ref_1543_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1543_index_offset_req_1;
      array_obj_ref_1543_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- unary operator type_cast_1492_inst
    process(add32_1483) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", add32_1483, tmp_var);
      type_cast_1492_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1506_inst
    process(shr_1503) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_1503, tmp_var);
      type_cast_1506_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1522_inst
    process(add76_1488) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", add76_1488, tmp_var);
      type_cast_1522_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1536_inst
    process(shr84_1533) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr84_1533, tmp_var);
      type_cast_1536_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1552_inst
    process(input_dim2x_x1_1478) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim2x_x1_1478, tmp_var);
      type_cast_1552_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1591_inst
    process(inc_1588) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_1588, tmp_var);
      type_cast_1591_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1617_inst
    process(inc109x_xinput_dim0x_x2_1607) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc109x_xinput_dim0x_x2_1607, tmp_var);
      type_cast_1617_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_1518_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1518_load_0_req_0;
      ptr_deref_1518_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1518_load_0_req_1;
      ptr_deref_1518_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1518_word_address_0;
      ptr_deref_1518_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_1547_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1547_store_0_req_0;
      ptr_deref_1547_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1547_store_0_req_1;
      ptr_deref_1547_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1547_word_address_0;
      data_in <= ptr_deref_1547_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block0_start_1326_inst RPIPE_Block0_start_1329_inst RPIPE_Block0_start_1347_inst RPIPE_Block0_start_1320_inst RPIPE_Block0_start_1317_inst RPIPE_Block0_start_1323_inst RPIPE_Block0_start_1332_inst RPIPE_Block0_start_1341_inst RPIPE_Block0_start_1335_inst RPIPE_Block0_start_1314_inst RPIPE_Block0_start_1344_inst RPIPE_Block0_start_1338_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(191 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 11 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 11 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 11 downto 0);
      signal guard_vector : std_logic_vector( 11 downto 0);
      constant outBUFs : IntegerArray(11 downto 0) := (11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(11 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false);
      constant guardBuffering: IntegerArray(11 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2);
      -- 
    begin -- 
      reqL_unguarded(11) <= RPIPE_Block0_start_1326_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block0_start_1329_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block0_start_1347_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block0_start_1320_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block0_start_1317_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block0_start_1323_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block0_start_1332_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block0_start_1341_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block0_start_1335_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block0_start_1314_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block0_start_1344_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block0_start_1338_inst_req_0;
      RPIPE_Block0_start_1326_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block0_start_1329_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block0_start_1347_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block0_start_1320_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block0_start_1317_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block0_start_1323_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block0_start_1332_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block0_start_1341_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block0_start_1335_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block0_start_1314_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block0_start_1344_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block0_start_1338_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(11) <= RPIPE_Block0_start_1326_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block0_start_1329_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block0_start_1347_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block0_start_1320_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block0_start_1317_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block0_start_1323_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block0_start_1332_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block0_start_1341_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block0_start_1335_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block0_start_1314_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block0_start_1344_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block0_start_1338_inst_req_1;
      RPIPE_Block0_start_1326_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block0_start_1329_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block0_start_1347_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block0_start_1320_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block0_start_1317_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block0_start_1323_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block0_start_1332_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block0_start_1341_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block0_start_1335_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block0_start_1314_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block0_start_1344_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block0_start_1338_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      call7_1327 <= data_out(191 downto 176);
      call9_1330 <= data_out(175 downto 160);
      call19_1348 <= data_out(159 downto 144);
      call3_1321 <= data_out(143 downto 128);
      call1_1318 <= data_out(127 downto 112);
      call5_1324 <= data_out(111 downto 96);
      call11_1333 <= data_out(95 downto 80);
      call15_1342 <= data_out(79 downto 64);
      call13_1336 <= data_out(63 downto 48);
      call_1315 <= data_out(47 downto 32);
      call17_1345 <= data_out(31 downto 16);
      call14_1339 <= data_out(15 downto 0);
      Block0_start_read_0_gI: SplitGuardInterface generic map(name => "Block0_start_read_0_gI", nreqs => 12, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_start_read_0: InputPortRevised -- 
        generic map ( name => "Block0_start_read_0", data_width => 16,  num_reqs => 12,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_start_pipe_read_req(0),
          oack => Block0_start_pipe_read_ack(0),
          odata => Block0_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block0_done_1633_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block0_done_1633_inst_req_0;
      WPIPE_Block0_done_1633_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block0_done_1633_inst_req_1;
      WPIPE_Block0_done_1633_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_1635_wire_constant;
      Block0_done_write_0_gI: SplitGuardInterface generic map(name => "Block0_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_done_pipe_write_req(0),
          oack => Block0_done_pipe_write_ack(0),
          odata => Block0_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeA_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeB is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeB;
architecture convTransposeB_arch of convTransposeB is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeB_CP_4133_start: Boolean;
  signal convTransposeB_CP_4133_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block1_start_1644_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1644_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1653_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1656_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1650_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1671_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1653_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1671_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1671_inst_req_0 : boolean;
  signal type_cast_1688_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1677_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1656_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1650_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1662_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1659_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1662_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1677_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1671_inst_req_1 : boolean;
  signal type_cast_1821_inst_ack_1 : boolean;
  signal type_cast_1696_inst_req_1 : boolean;
  signal type_cast_1696_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1647_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1659_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1665_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1668_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1668_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1656_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1665_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1656_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1653_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1647_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1644_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1653_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1665_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1665_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1659_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1647_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1644_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1662_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1662_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1647_inst_ack_1 : boolean;
  signal type_cast_1692_inst_req_0 : boolean;
  signal type_cast_1692_inst_ack_0 : boolean;
  signal type_cast_1692_inst_ack_1 : boolean;
  signal type_cast_1821_inst_req_0 : boolean;
  signal type_cast_1821_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1668_inst_ack_1 : boolean;
  signal type_cast_1835_inst_req_1 : boolean;
  signal type_cast_1835_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1668_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1650_inst_ack_0 : boolean;
  signal type_cast_1835_inst_req_0 : boolean;
  signal type_cast_1835_inst_ack_0 : boolean;
  signal type_cast_1692_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1674_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1659_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1674_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1650_inst_req_0 : boolean;
  signal type_cast_1696_inst_req_0 : boolean;
  signal type_cast_1696_inst_ack_0 : boolean;
  signal type_cast_1821_inst_req_1 : boolean;
  signal type_cast_1688_inst_ack_0 : boolean;
  signal type_cast_1688_inst_ack_1 : boolean;
  signal type_cast_1688_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1674_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1674_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1677_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1677_inst_req_0 : boolean;
  signal array_obj_ref_1841_index_offset_req_0 : boolean;
  signal array_obj_ref_1841_index_offset_ack_0 : boolean;
  signal array_obj_ref_1841_index_offset_req_1 : boolean;
  signal array_obj_ref_1841_index_offset_ack_1 : boolean;
  signal addr_of_1842_final_reg_req_0 : boolean;
  signal addr_of_1842_final_reg_ack_0 : boolean;
  signal addr_of_1842_final_reg_req_1 : boolean;
  signal addr_of_1842_final_reg_ack_1 : boolean;
  signal ptr_deref_1846_load_0_req_0 : boolean;
  signal ptr_deref_1846_load_0_ack_0 : boolean;
  signal ptr_deref_1846_load_0_req_1 : boolean;
  signal ptr_deref_1846_load_0_ack_1 : boolean;
  signal type_cast_1851_inst_req_0 : boolean;
  signal type_cast_1851_inst_ack_0 : boolean;
  signal type_cast_1851_inst_req_1 : boolean;
  signal type_cast_1851_inst_ack_1 : boolean;
  signal type_cast_1865_inst_req_0 : boolean;
  signal type_cast_1865_inst_ack_0 : boolean;
  signal type_cast_1865_inst_req_1 : boolean;
  signal type_cast_1865_inst_ack_1 : boolean;
  signal array_obj_ref_1871_index_offset_req_0 : boolean;
  signal array_obj_ref_1871_index_offset_ack_0 : boolean;
  signal array_obj_ref_1871_index_offset_req_1 : boolean;
  signal array_obj_ref_1871_index_offset_ack_1 : boolean;
  signal addr_of_1872_final_reg_req_0 : boolean;
  signal addr_of_1872_final_reg_ack_0 : boolean;
  signal addr_of_1872_final_reg_req_1 : boolean;
  signal addr_of_1872_final_reg_ack_1 : boolean;
  signal ptr_deref_1875_store_0_req_0 : boolean;
  signal ptr_deref_1875_store_0_ack_0 : boolean;
  signal ptr_deref_1875_store_0_req_1 : boolean;
  signal ptr_deref_1875_store_0_ack_1 : boolean;
  signal type_cast_1881_inst_req_0 : boolean;
  signal type_cast_1881_inst_ack_0 : boolean;
  signal type_cast_1881_inst_req_1 : boolean;
  signal type_cast_1881_inst_ack_1 : boolean;
  signal if_stmt_1896_branch_req_0 : boolean;
  signal if_stmt_1896_branch_ack_1 : boolean;
  signal if_stmt_1896_branch_ack_0 : boolean;
  signal type_cast_1920_inst_req_0 : boolean;
  signal type_cast_1920_inst_ack_0 : boolean;
  signal type_cast_1920_inst_req_1 : boolean;
  signal type_cast_1920_inst_ack_1 : boolean;
  signal type_cast_1935_inst_req_0 : boolean;
  signal type_cast_1935_inst_ack_0 : boolean;
  signal type_cast_1935_inst_req_1 : boolean;
  signal type_cast_1935_inst_ack_1 : boolean;
  signal type_cast_1945_inst_req_0 : boolean;
  signal type_cast_1945_inst_ack_0 : boolean;
  signal type_cast_1945_inst_req_1 : boolean;
  signal type_cast_1945_inst_ack_1 : boolean;
  signal if_stmt_1952_branch_req_0 : boolean;
  signal if_stmt_1952_branch_ack_1 : boolean;
  signal if_stmt_1952_branch_ack_0 : boolean;
  signal WPIPE_Block1_done_1960_inst_req_0 : boolean;
  signal WPIPE_Block1_done_1960_inst_ack_0 : boolean;
  signal WPIPE_Block1_done_1960_inst_req_1 : boolean;
  signal WPIPE_Block1_done_1960_inst_ack_1 : boolean;
  signal type_cast_1731_inst_req_0 : boolean;
  signal type_cast_1731_inst_ack_0 : boolean;
  signal type_cast_1731_inst_req_1 : boolean;
  signal type_cast_1731_inst_ack_1 : boolean;
  signal phi_stmt_1728_req_0 : boolean;
  signal phi_stmt_1734_req_0 : boolean;
  signal type_cast_1733_inst_req_0 : boolean;
  signal type_cast_1733_inst_ack_0 : boolean;
  signal type_cast_1733_inst_req_1 : boolean;
  signal type_cast_1733_inst_ack_1 : boolean;
  signal phi_stmt_1728_req_1 : boolean;
  signal type_cast_1740_inst_req_0 : boolean;
  signal type_cast_1740_inst_ack_0 : boolean;
  signal type_cast_1740_inst_req_1 : boolean;
  signal type_cast_1740_inst_ack_1 : boolean;
  signal phi_stmt_1734_req_1 : boolean;
  signal phi_stmt_1728_ack_0 : boolean;
  signal phi_stmt_1734_ack_0 : boolean;
  signal type_cast_1797_inst_req_0 : boolean;
  signal type_cast_1797_inst_ack_0 : boolean;
  signal type_cast_1797_inst_req_1 : boolean;
  signal type_cast_1797_inst_ack_1 : boolean;
  signal phi_stmt_1794_req_0 : boolean;
  signal phi_stmt_1794_req_1 : boolean;
  signal phi_stmt_1794_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeB_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeB_CP_4133_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeB_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_4133_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeB_CP_4133_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_4133_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeB_CP_4133: Block -- control-path 
    signal convTransposeB_CP_4133_elements: BooleanArray(89 downto 0);
    -- 
  begin -- 
    convTransposeB_CP_4133_elements(0) <= convTransposeB_CP_4133_start;
    convTransposeB_CP_4133_symbol <= convTransposeB_CP_4133_elements(67);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1644_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1644_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1644_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1642/$entry
      -- CP-element group 0: 	 branch_block_stmt_1642/branch_block_stmt_1642__entry__
      -- CP-element group 0: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678__entry__
      -- 
    rr_4181_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4181_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(0), ack => RPIPE_Block1_start_1644_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1644_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1644_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1644_update_start_
      -- CP-element group 1: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1644_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1644_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1644_sample_completed_
      -- 
    ra_4182_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1644_inst_ack_0, ack => convTransposeB_CP_4133_elements(1)); -- 
    cr_4186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(1), ack => RPIPE_Block1_start_1644_inst_req_1); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1644_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1644_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1644_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1647_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1647_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1647_sample_start_
      -- 
    ca_4187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1644_inst_ack_1, ack => convTransposeB_CP_4133_elements(2)); -- 
    rr_4195_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4195_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(2), ack => RPIPE_Block1_start_1647_inst_req_0); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1647_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1647_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1647_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1647_Update/cr
      -- CP-element group 3: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1647_update_start_
      -- CP-element group 3: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1647_sample_completed_
      -- 
    ra_4196_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1647_inst_ack_0, ack => convTransposeB_CP_4133_elements(3)); -- 
    cr_4200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(3), ack => RPIPE_Block1_start_1647_inst_req_1); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1650_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1650_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1647_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1647_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1650_Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1647_update_completed_
      -- 
    ca_4201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1647_inst_ack_1, ack => convTransposeB_CP_4133_elements(4)); -- 
    rr_4209_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4209_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(4), ack => RPIPE_Block1_start_1650_inst_req_0); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1650_Update/cr
      -- CP-element group 5: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1650_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1650_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1650_update_start_
      -- CP-element group 5: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1650_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1650_Sample/ra
      -- 
    ra_4210_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1650_inst_ack_0, ack => convTransposeB_CP_4133_elements(5)); -- 
    cr_4214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(5), ack => RPIPE_Block1_start_1650_inst_req_1); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1650_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1653_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1653_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1653_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1650_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1650_update_completed_
      -- 
    ca_4215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1650_inst_ack_1, ack => convTransposeB_CP_4133_elements(6)); -- 
    rr_4223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(6), ack => RPIPE_Block1_start_1653_inst_req_0); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1653_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1653_Sample/ra
      -- CP-element group 7: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1653_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1653_Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1653_update_start_
      -- CP-element group 7: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1653_Update/cr
      -- 
    ra_4224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1653_inst_ack_0, ack => convTransposeB_CP_4133_elements(7)); -- 
    cr_4228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(7), ack => RPIPE_Block1_start_1653_inst_req_1); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1656_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1653_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1653_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1656_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1653_Update/ca
      -- CP-element group 8: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1656_sample_start_
      -- 
    ca_4229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1653_inst_ack_1, ack => convTransposeB_CP_4133_elements(8)); -- 
    rr_4237_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4237_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(8), ack => RPIPE_Block1_start_1656_inst_req_0); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1656_update_start_
      -- CP-element group 9: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1656_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1656_Update/cr
      -- CP-element group 9: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1656_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1656_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1656_sample_completed_
      -- 
    ra_4238_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1656_inst_ack_0, ack => convTransposeB_CP_4133_elements(9)); -- 
    cr_4242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(9), ack => RPIPE_Block1_start_1656_inst_req_1); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1656_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1656_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1659_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1656_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1659_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1659_Sample/rr
      -- 
    ca_4243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1656_inst_ack_1, ack => convTransposeB_CP_4133_elements(10)); -- 
    rr_4251_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4251_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(10), ack => RPIPE_Block1_start_1659_inst_req_0); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1659_Update/cr
      -- CP-element group 11: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1659_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1659_update_start_
      -- CP-element group 11: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1659_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1659_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1659_Sample/ra
      -- 
    ra_4252_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1659_inst_ack_0, ack => convTransposeB_CP_4133_elements(11)); -- 
    cr_4256_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4256_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(11), ack => RPIPE_Block1_start_1659_inst_req_1); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1659_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1662_sample_start_
      -- CP-element group 12: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1659_Update/ca
      -- CP-element group 12: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1659_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1662_Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1662_Sample/rr
      -- 
    ca_4257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1659_inst_ack_1, ack => convTransposeB_CP_4133_elements(12)); -- 
    rr_4265_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4265_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(12), ack => RPIPE_Block1_start_1662_inst_req_0); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1662_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1662_update_start_
      -- CP-element group 13: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1662_Update/cr
      -- CP-element group 13: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1662_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1662_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1662_Sample/ra
      -- 
    ra_4266_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1662_inst_ack_0, ack => convTransposeB_CP_4133_elements(13)); -- 
    cr_4270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(13), ack => RPIPE_Block1_start_1662_inst_req_1); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1665_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1662_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1665_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1662_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1665_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1662_Update/$exit
      -- 
    ca_4271_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1662_inst_ack_1, ack => convTransposeB_CP_4133_elements(14)); -- 
    rr_4279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(14), ack => RPIPE_Block1_start_1665_inst_req_0); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1665_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1665_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1665_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1665_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1665_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1665_Update/$entry
      -- 
    ra_4280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1665_inst_ack_0, ack => convTransposeB_CP_4133_elements(15)); -- 
    cr_4284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(15), ack => RPIPE_Block1_start_1665_inst_req_1); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1665_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1668_Sample/$entry
      -- CP-element group 16: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1668_Sample/rr
      -- CP-element group 16: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1665_Update/ca
      -- CP-element group 16: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1668_sample_start_
      -- CP-element group 16: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1665_Update/$exit
      -- 
    ca_4285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1665_inst_ack_1, ack => convTransposeB_CP_4133_elements(16)); -- 
    rr_4293_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4293_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(16), ack => RPIPE_Block1_start_1668_inst_req_0); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1668_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1668_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1668_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1668_update_start_
      -- CP-element group 17: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1668_Update/cr
      -- CP-element group 17: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1668_Update/$entry
      -- 
    ra_4294_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1668_inst_ack_0, ack => convTransposeB_CP_4133_elements(17)); -- 
    cr_4298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(17), ack => RPIPE_Block1_start_1668_inst_req_1); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1671_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1671_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1668_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1671_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1668_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1668_Update/$exit
      -- 
    ca_4299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1668_inst_ack_1, ack => convTransposeB_CP_4133_elements(18)); -- 
    rr_4307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(18), ack => RPIPE_Block1_start_1671_inst_req_0); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1671_Update/$entry
      -- CP-element group 19: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1671_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1671_Sample/ra
      -- CP-element group 19: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1671_Update/cr
      -- CP-element group 19: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1671_update_start_
      -- CP-element group 19: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1671_sample_completed_
      -- 
    ra_4308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1671_inst_ack_0, ack => convTransposeB_CP_4133_elements(19)); -- 
    cr_4312_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4312_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(19), ack => RPIPE_Block1_start_1671_inst_req_1); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1674_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1671_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1671_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1674_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1671_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1674_Sample/rr
      -- 
    ca_4313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1671_inst_ack_1, ack => convTransposeB_CP_4133_elements(20)); -- 
    rr_4321_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4321_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(20), ack => RPIPE_Block1_start_1674_inst_req_0); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1674_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1674_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1674_update_start_
      -- CP-element group 21: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1674_Update/cr
      -- CP-element group 21: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1674_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1674_Sample/ra
      -- 
    ra_4322_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1674_inst_ack_0, ack => convTransposeB_CP_4133_elements(21)); -- 
    cr_4326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(21), ack => RPIPE_Block1_start_1674_inst_req_1); -- 
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (6) 
      -- CP-element group 22: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1674_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1677_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1677_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1674_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1674_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1677_Sample/rr
      -- 
    ca_4327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1674_inst_ack_1, ack => convTransposeB_CP_4133_elements(22)); -- 
    rr_4335_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4335_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(22), ack => RPIPE_Block1_start_1677_inst_req_0); -- 
    -- CP-element group 23:  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (6) 
      -- CP-element group 23: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1677_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1677_Update/cr
      -- CP-element group 23: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1677_update_start_
      -- CP-element group 23: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1677_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1677_Update/$entry
      -- CP-element group 23: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1677_Sample/ra
      -- 
    ra_4336_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1677_inst_ack_0, ack => convTransposeB_CP_4133_elements(23)); -- 
    cr_4340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(23), ack => RPIPE_Block1_start_1677_inst_req_1); -- 
    -- CP-element group 24:  fork  transition  place  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24: 	26 
    -- CP-element group 24: 	27 
    -- CP-element group 24: 	28 
    -- CP-element group 24: 	29 
    -- CP-element group 24: 	30 
    -- CP-element group 24:  members (25) 
      -- CP-element group 24: 	 branch_block_stmt_1642/assign_stmt_1685_to_assign_stmt_1725/$entry
      -- CP-element group 24: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1677_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_1642/assign_stmt_1685_to_assign_stmt_1725/type_cast_1696_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1642/assign_stmt_1685_to_assign_stmt_1725/type_cast_1688_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1677_Update/ca
      -- CP-element group 24: 	 branch_block_stmt_1642/assign_stmt_1685_to_assign_stmt_1725/type_cast_1692_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1642/assign_stmt_1685_to_assign_stmt_1725/type_cast_1696_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_1642/assign_stmt_1685_to_assign_stmt_1725/type_cast_1692_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1642/assign_stmt_1685_to_assign_stmt_1725/type_cast_1692_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_1642/assign_stmt_1685_to_assign_stmt_1725/type_cast_1688_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1642/assign_stmt_1685_to_assign_stmt_1725/type_cast_1692_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1642/assign_stmt_1685_to_assign_stmt_1725/type_cast_1692_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_1642/assign_stmt_1685_to_assign_stmt_1725/type_cast_1696_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1642/assign_stmt_1685_to_assign_stmt_1725/type_cast_1696_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_1642/assign_stmt_1685_to_assign_stmt_1725/type_cast_1696_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1642/assign_stmt_1685_to_assign_stmt_1725/type_cast_1692_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_1642/assign_stmt_1685_to_assign_stmt_1725/type_cast_1696_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_1642/assign_stmt_1685_to_assign_stmt_1725/type_cast_1688_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1642/assign_stmt_1685_to_assign_stmt_1725/type_cast_1688_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_1642/assign_stmt_1685_to_assign_stmt_1725/type_cast_1688_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1642/assign_stmt_1685_to_assign_stmt_1725/type_cast_1688_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/RPIPE_Block1_start_1677_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678/$exit
      -- CP-element group 24: 	 branch_block_stmt_1642/assign_stmt_1645_to_assign_stmt_1678__exit__
      -- CP-element group 24: 	 branch_block_stmt_1642/assign_stmt_1685_to_assign_stmt_1725__entry__
      -- 
    ca_4341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1677_inst_ack_1, ack => convTransposeB_CP_4133_elements(24)); -- 
    rr_4352_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4352_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(24), ack => type_cast_1688_inst_req_0); -- 
    cr_4385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(24), ack => type_cast_1696_inst_req_1); -- 
    rr_4366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(24), ack => type_cast_1692_inst_req_0); -- 
    cr_4371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(24), ack => type_cast_1692_inst_req_1); -- 
    rr_4380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(24), ack => type_cast_1696_inst_req_0); -- 
    cr_4357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(24), ack => type_cast_1688_inst_req_1); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_1642/assign_stmt_1685_to_assign_stmt_1725/type_cast_1688_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_1642/assign_stmt_1685_to_assign_stmt_1725/type_cast_1688_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_1642/assign_stmt_1685_to_assign_stmt_1725/type_cast_1688_Sample/ra
      -- 
    ra_4353_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1688_inst_ack_0, ack => convTransposeB_CP_4133_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	31 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1642/assign_stmt_1685_to_assign_stmt_1725/type_cast_1688_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_1642/assign_stmt_1685_to_assign_stmt_1725/type_cast_1688_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_1642/assign_stmt_1685_to_assign_stmt_1725/type_cast_1688_Update/ca
      -- 
    ca_4358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1688_inst_ack_1, ack => convTransposeB_CP_4133_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	24 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1642/assign_stmt_1685_to_assign_stmt_1725/type_cast_1692_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_1642/assign_stmt_1685_to_assign_stmt_1725/type_cast_1692_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_1642/assign_stmt_1685_to_assign_stmt_1725/type_cast_1692_Sample/ra
      -- 
    ra_4367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1692_inst_ack_0, ack => convTransposeB_CP_4133_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	24 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	31 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1642/assign_stmt_1685_to_assign_stmt_1725/type_cast_1692_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_1642/assign_stmt_1685_to_assign_stmt_1725/type_cast_1692_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_1642/assign_stmt_1685_to_assign_stmt_1725/type_cast_1692_Update/ca
      -- 
    ca_4372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1692_inst_ack_1, ack => convTransposeB_CP_4133_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	24 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_1642/assign_stmt_1685_to_assign_stmt_1725/type_cast_1696_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_1642/assign_stmt_1685_to_assign_stmt_1725/type_cast_1696_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_1642/assign_stmt_1685_to_assign_stmt_1725/type_cast_1696_Sample/ra
      -- 
    ra_4381_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1696_inst_ack_0, ack => convTransposeB_CP_4133_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	24 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1642/assign_stmt_1685_to_assign_stmt_1725/type_cast_1696_Update/ca
      -- CP-element group 30: 	 branch_block_stmt_1642/assign_stmt_1685_to_assign_stmt_1725/type_cast_1696_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_1642/assign_stmt_1685_to_assign_stmt_1725/type_cast_1696_Update/$exit
      -- 
    ca_4386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1696_inst_ack_1, ack => convTransposeB_CP_4133_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  place  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	26 
    -- CP-element group 31: 	28 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	68 
    -- CP-element group 31: 	69 
    -- CP-element group 31: 	71 
    -- CP-element group 31:  members (14) 
      -- CP-element group 31: 	 branch_block_stmt_1642/assign_stmt_1685_to_assign_stmt_1725/$exit
      -- CP-element group 31: 	 branch_block_stmt_1642/assign_stmt_1685_to_assign_stmt_1725__exit__
      -- CP-element group 31: 	 branch_block_stmt_1642/entry_whilex_xbodyx_xouter
      -- CP-element group 31: 	 branch_block_stmt_1642/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 31: 	 branch_block_stmt_1642/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1728/$entry
      -- CP-element group 31: 	 branch_block_stmt_1642/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/$entry
      -- CP-element group 31: 	 branch_block_stmt_1642/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1731/$entry
      -- CP-element group 31: 	 branch_block_stmt_1642/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1731/SplitProtocol/$entry
      -- CP-element group 31: 	 branch_block_stmt_1642/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1731/SplitProtocol/Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1642/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1731/SplitProtocol/Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_1642/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1731/SplitProtocol/Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_1642/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1731/SplitProtocol/Update/cr
      -- CP-element group 31: 	 branch_block_stmt_1642/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/$entry
      -- CP-element group 31: 	 branch_block_stmt_1642/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/$entry
      -- 
    rr_4776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(31), ack => type_cast_1731_inst_req_0); -- 
    cr_4781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(31), ack => type_cast_1731_inst_req_1); -- 
    convTransposeB_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4133_elements(26) & convTransposeB_CP_4133_elements(28) & convTransposeB_CP_4133_elements(30);
      gj_convTransposeB_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4133_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	89 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1821_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1821_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1821_sample_completed_
      -- 
    ra_4401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1821_inst_ack_0, ack => convTransposeB_CP_4133_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	89 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1821_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1821_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1835_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1821_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1835_Sample/rr
      -- CP-element group 33: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1835_sample_start_
      -- 
    ca_4406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1821_inst_ack_1, ack => convTransposeB_CP_4133_elements(33)); -- 
    rr_4414_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4414_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(33), ack => type_cast_1835_inst_req_0); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1835_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1835_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1835_Sample/ra
      -- 
    ra_4415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1835_inst_ack_0, ack => convTransposeB_CP_4133_elements(34)); -- 
    -- CP-element group 35:  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	89 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (16) 
      -- CP-element group 35: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1835_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1841_index_computed_1
      -- CP-element group 35: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1841_index_resized_1
      -- CP-element group 35: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1841_index_scaled_1
      -- CP-element group 35: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1841_index_resize_1/index_resize_req
      -- CP-element group 35: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1841_index_resize_1/index_resize_ack
      -- CP-element group 35: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1835_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1835_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1841_index_resize_1/$entry
      -- CP-element group 35: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1841_index_resize_1/$exit
      -- CP-element group 35: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1841_index_scale_1/$entry
      -- CP-element group 35: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1841_index_scale_1/$exit
      -- CP-element group 35: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1841_index_scale_1/scale_rename_req
      -- CP-element group 35: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1841_index_scale_1/scale_rename_ack
      -- CP-element group 35: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1841_final_index_sum_regn_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1841_final_index_sum_regn_Sample/req
      -- 
    ca_4420_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1835_inst_ack_1, ack => convTransposeB_CP_4133_elements(35)); -- 
    req_4445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(35), ack => array_obj_ref_1841_index_offset_req_0); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	55 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1841_final_index_sum_regn_sample_complete
      -- CP-element group 36: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1841_final_index_sum_regn_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1841_final_index_sum_regn_Sample/ack
      -- 
    ack_4446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1841_index_offset_ack_0, ack => convTransposeB_CP_4133_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	89 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (11) 
      -- CP-element group 37: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/addr_of_1842_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1841_root_address_calculated
      -- CP-element group 37: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1841_offset_calculated
      -- CP-element group 37: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1841_final_index_sum_regn_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1841_final_index_sum_regn_Update/ack
      -- CP-element group 37: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1841_base_plus_offset/$entry
      -- CP-element group 37: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1841_base_plus_offset/$exit
      -- CP-element group 37: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1841_base_plus_offset/sum_rename_req
      -- CP-element group 37: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1841_base_plus_offset/sum_rename_ack
      -- CP-element group 37: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/addr_of_1842_request/$entry
      -- CP-element group 37: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/addr_of_1842_request/req
      -- 
    ack_4451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1841_index_offset_ack_1, ack => convTransposeB_CP_4133_elements(37)); -- 
    req_4460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(37), ack => addr_of_1842_final_reg_req_0); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/addr_of_1842_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/addr_of_1842_request/$exit
      -- CP-element group 38: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/addr_of_1842_request/ack
      -- 
    ack_4461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1842_final_reg_ack_0, ack => convTransposeB_CP_4133_elements(38)); -- 
    -- CP-element group 39:  join  fork  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	89 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (24) 
      -- CP-element group 39: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/addr_of_1842_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/addr_of_1842_complete/$exit
      -- CP-element group 39: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/addr_of_1842_complete/ack
      -- CP-element group 39: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1846_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1846_base_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1846_word_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1846_root_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1846_base_address_resized
      -- CP-element group 39: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1846_base_addr_resize/$entry
      -- CP-element group 39: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1846_base_addr_resize/$exit
      -- CP-element group 39: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1846_base_addr_resize/base_resize_req
      -- CP-element group 39: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1846_base_addr_resize/base_resize_ack
      -- CP-element group 39: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1846_base_plus_offset/$entry
      -- CP-element group 39: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1846_base_plus_offset/$exit
      -- CP-element group 39: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1846_base_plus_offset/sum_rename_req
      -- CP-element group 39: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1846_base_plus_offset/sum_rename_ack
      -- CP-element group 39: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1846_word_addrgen/$entry
      -- CP-element group 39: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1846_word_addrgen/$exit
      -- CP-element group 39: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1846_word_addrgen/root_register_req
      -- CP-element group 39: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1846_word_addrgen/root_register_ack
      -- CP-element group 39: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1846_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1846_Sample/word_access_start/$entry
      -- CP-element group 39: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1846_Sample/word_access_start/word_0/$entry
      -- CP-element group 39: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1846_Sample/word_access_start/word_0/rr
      -- 
    ack_4466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1842_final_reg_ack_1, ack => convTransposeB_CP_4133_elements(39)); -- 
    rr_4499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(39), ack => ptr_deref_1846_load_0_req_0); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (5) 
      -- CP-element group 40: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1846_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1846_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1846_Sample/word_access_start/$exit
      -- CP-element group 40: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1846_Sample/word_access_start/word_0/$exit
      -- CP-element group 40: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1846_Sample/word_access_start/word_0/ra
      -- 
    ra_4500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1846_load_0_ack_0, ack => convTransposeB_CP_4133_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	89 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	50 
    -- CP-element group 41:  members (9) 
      -- CP-element group 41: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1846_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1846_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1846_Update/word_access_complete/$exit
      -- CP-element group 41: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1846_Update/word_access_complete/word_0/$exit
      -- CP-element group 41: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1846_Update/word_access_complete/word_0/ca
      -- CP-element group 41: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1846_Update/ptr_deref_1846_Merge/$entry
      -- CP-element group 41: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1846_Update/ptr_deref_1846_Merge/$exit
      -- CP-element group 41: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1846_Update/ptr_deref_1846_Merge/merge_req
      -- CP-element group 41: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1846_Update/ptr_deref_1846_Merge/merge_ack
      -- 
    ca_4511_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1846_load_0_ack_1, ack => convTransposeB_CP_4133_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	89 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1851_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1851_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1851_Sample/ra
      -- 
    ra_4525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1851_inst_ack_0, ack => convTransposeB_CP_4133_elements(42)); -- 
    -- CP-element group 43:  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	89 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (6) 
      -- CP-element group 43: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1851_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1851_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1851_Update/ca
      -- CP-element group 43: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1865_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1865_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1865_Sample/rr
      -- 
    ca_4530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1851_inst_ack_1, ack => convTransposeB_CP_4133_elements(43)); -- 
    rr_4538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(43), ack => type_cast_1865_inst_req_0); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1865_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1865_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1865_Sample/ra
      -- 
    ra_4539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1865_inst_ack_0, ack => convTransposeB_CP_4133_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	89 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (16) 
      -- CP-element group 45: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1871_index_scale_1/$entry
      -- CP-element group 45: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1865_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1865_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1865_Update/ca
      -- CP-element group 45: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1871_index_resized_1
      -- CP-element group 45: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1871_index_scaled_1
      -- CP-element group 45: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1871_index_computed_1
      -- CP-element group 45: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1871_index_resize_1/$entry
      -- CP-element group 45: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1871_index_resize_1/$exit
      -- CP-element group 45: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1871_index_resize_1/index_resize_req
      -- CP-element group 45: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1871_index_resize_1/index_resize_ack
      -- CP-element group 45: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1871_index_scale_1/$exit
      -- CP-element group 45: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1871_index_scale_1/scale_rename_req
      -- CP-element group 45: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1871_index_scale_1/scale_rename_ack
      -- CP-element group 45: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1871_final_index_sum_regn_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1871_final_index_sum_regn_Sample/req
      -- 
    ca_4544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1865_inst_ack_1, ack => convTransposeB_CP_4133_elements(45)); -- 
    req_4569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(45), ack => array_obj_ref_1871_index_offset_req_0); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	55 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1871_final_index_sum_regn_sample_complete
      -- CP-element group 46: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1871_final_index_sum_regn_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1871_final_index_sum_regn_Sample/ack
      -- 
    ack_4570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1871_index_offset_ack_0, ack => convTransposeB_CP_4133_elements(46)); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	89 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (11) 
      -- CP-element group 47: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/addr_of_1872_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1871_root_address_calculated
      -- CP-element group 47: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1871_offset_calculated
      -- CP-element group 47: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1871_final_index_sum_regn_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1871_final_index_sum_regn_Update/ack
      -- CP-element group 47: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1871_base_plus_offset/$entry
      -- CP-element group 47: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1871_base_plus_offset/$exit
      -- CP-element group 47: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1871_base_plus_offset/sum_rename_req
      -- CP-element group 47: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1871_base_plus_offset/sum_rename_ack
      -- CP-element group 47: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/addr_of_1872_request/$entry
      -- CP-element group 47: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/addr_of_1872_request/req
      -- 
    ack_4575_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1871_index_offset_ack_1, ack => convTransposeB_CP_4133_elements(47)); -- 
    req_4584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(47), ack => addr_of_1872_final_reg_req_0); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/addr_of_1872_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/addr_of_1872_request/$exit
      -- CP-element group 48: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/addr_of_1872_request/ack
      -- 
    ack_4585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1872_final_reg_ack_0, ack => convTransposeB_CP_4133_elements(48)); -- 
    -- CP-element group 49:  fork  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	89 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (19) 
      -- CP-element group 49: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/addr_of_1872_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/addr_of_1872_complete/$exit
      -- CP-element group 49: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/addr_of_1872_complete/ack
      -- CP-element group 49: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1875_base_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1875_word_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1875_root_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1875_base_address_resized
      -- CP-element group 49: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1875_base_addr_resize/$entry
      -- CP-element group 49: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1875_base_addr_resize/$exit
      -- CP-element group 49: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1875_base_addr_resize/base_resize_req
      -- CP-element group 49: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1875_base_addr_resize/base_resize_ack
      -- CP-element group 49: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1875_base_plus_offset/$entry
      -- CP-element group 49: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1875_base_plus_offset/$exit
      -- CP-element group 49: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1875_base_plus_offset/sum_rename_req
      -- CP-element group 49: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1875_base_plus_offset/sum_rename_ack
      -- CP-element group 49: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1875_word_addrgen/$entry
      -- CP-element group 49: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1875_word_addrgen/$exit
      -- CP-element group 49: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1875_word_addrgen/root_register_req
      -- CP-element group 49: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1875_word_addrgen/root_register_ack
      -- 
    ack_4590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1872_final_reg_ack_1, ack => convTransposeB_CP_4133_elements(49)); -- 
    -- CP-element group 50:  join  transition  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	41 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1875_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1875_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1875_Sample/ptr_deref_1875_Split/$entry
      -- CP-element group 50: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1875_Sample/ptr_deref_1875_Split/$exit
      -- CP-element group 50: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1875_Sample/ptr_deref_1875_Split/split_req
      -- CP-element group 50: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1875_Sample/ptr_deref_1875_Split/split_ack
      -- CP-element group 50: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1875_Sample/word_access_start/$entry
      -- CP-element group 50: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1875_Sample/word_access_start/word_0/$entry
      -- CP-element group 50: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1875_Sample/word_access_start/word_0/rr
      -- 
    rr_4628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(50), ack => ptr_deref_1875_store_0_req_0); -- 
    convTransposeB_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4133_elements(41) & convTransposeB_CP_4133_elements(49);
      gj_convTransposeB_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4133_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (5) 
      -- CP-element group 51: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1875_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1875_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1875_Sample/word_access_start/$exit
      -- CP-element group 51: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1875_Sample/word_access_start/word_0/$exit
      -- CP-element group 51: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1875_Sample/word_access_start/word_0/ra
      -- 
    ra_4629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1875_store_0_ack_0, ack => convTransposeB_CP_4133_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	89 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	55 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1875_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1875_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1875_Update/word_access_complete/$exit
      -- CP-element group 52: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1875_Update/word_access_complete/word_0/$exit
      -- CP-element group 52: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1875_Update/word_access_complete/word_0/ca
      -- 
    ca_4640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1875_store_0_ack_1, ack => convTransposeB_CP_4133_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	89 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1881_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1881_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1881_Sample/ra
      -- 
    ra_4649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1881_inst_ack_0, ack => convTransposeB_CP_4133_elements(53)); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	89 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1881_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1881_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1881_Update/ca
      -- 
    ca_4654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1881_inst_ack_1, ack => convTransposeB_CP_4133_elements(54)); -- 
    -- CP-element group 55:  branch  join  transition  place  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	36 
    -- CP-element group 55: 	46 
    -- CP-element group 55: 	52 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (10) 
      -- CP-element group 55: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/$exit
      -- CP-element group 55: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895__exit__
      -- CP-element group 55: 	 branch_block_stmt_1642/if_stmt_1896__entry__
      -- CP-element group 55: 	 branch_block_stmt_1642/if_stmt_1896_dead_link/$entry
      -- CP-element group 55: 	 branch_block_stmt_1642/if_stmt_1896_eval_test/$entry
      -- CP-element group 55: 	 branch_block_stmt_1642/if_stmt_1896_eval_test/$exit
      -- CP-element group 55: 	 branch_block_stmt_1642/if_stmt_1896_eval_test/branch_req
      -- CP-element group 55: 	 branch_block_stmt_1642/R_cmp_1897_place
      -- CP-element group 55: 	 branch_block_stmt_1642/if_stmt_1896_if_link/$entry
      -- CP-element group 55: 	 branch_block_stmt_1642/if_stmt_1896_else_link/$entry
      -- 
    branch_req_4662_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4662_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(55), ack => if_stmt_1896_branch_req_0); -- 
    convTransposeB_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4133_elements(36) & convTransposeB_CP_4133_elements(46) & convTransposeB_CP_4133_elements(52) & convTransposeB_CP_4133_elements(54);
      gj_convTransposeB_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4133_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	84 
    -- CP-element group 56: 	85 
    -- CP-element group 56:  members (24) 
      -- CP-element group 56: 	 branch_block_stmt_1642/merge_stmt_1902__exit__
      -- CP-element group 56: 	 branch_block_stmt_1642/assign_stmt_1908__entry__
      -- CP-element group 56: 	 branch_block_stmt_1642/assign_stmt_1908__exit__
      -- CP-element group 56: 	 branch_block_stmt_1642/ifx_xthen_whilex_xbody
      -- CP-element group 56: 	 branch_block_stmt_1642/if_stmt_1896_if_link/$exit
      -- CP-element group 56: 	 branch_block_stmt_1642/if_stmt_1896_if_link/if_choice_transition
      -- CP-element group 56: 	 branch_block_stmt_1642/whilex_xbody_ifx_xthen
      -- CP-element group 56: 	 branch_block_stmt_1642/assign_stmt_1908/$entry
      -- CP-element group 56: 	 branch_block_stmt_1642/assign_stmt_1908/$exit
      -- CP-element group 56: 	 branch_block_stmt_1642/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 56: 	 branch_block_stmt_1642/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1794/$entry
      -- CP-element group 56: 	 branch_block_stmt_1642/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/$entry
      -- CP-element group 56: 	 branch_block_stmt_1642/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/type_cast_1797/$entry
      -- CP-element group 56: 	 branch_block_stmt_1642/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/type_cast_1797/SplitProtocol/$entry
      -- CP-element group 56: 	 branch_block_stmt_1642/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/type_cast_1797/SplitProtocol/Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_1642/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/type_cast_1797/SplitProtocol/Sample/rr
      -- CP-element group 56: 	 branch_block_stmt_1642/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/type_cast_1797/SplitProtocol/Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_1642/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/type_cast_1797/SplitProtocol/Update/cr
      -- CP-element group 56: 	 branch_block_stmt_1642/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 56: 	 branch_block_stmt_1642/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 56: 	 branch_block_stmt_1642/merge_stmt_1902_PhiReqMerge
      -- CP-element group 56: 	 branch_block_stmt_1642/merge_stmt_1902_PhiAck/$entry
      -- CP-element group 56: 	 branch_block_stmt_1642/merge_stmt_1902_PhiAck/$exit
      -- CP-element group 56: 	 branch_block_stmt_1642/merge_stmt_1902_PhiAck/dummy
      -- 
    if_choice_transition_4667_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1896_branch_ack_1, ack => convTransposeB_CP_4133_elements(56)); -- 
    rr_4865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(56), ack => type_cast_1797_inst_req_0); -- 
    cr_4870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(56), ack => type_cast_1797_inst_req_1); -- 
    -- CP-element group 57:  fork  transition  place  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57: 	59 
    -- CP-element group 57: 	61 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (24) 
      -- CP-element group 57: 	 branch_block_stmt_1642/merge_stmt_1910__exit__
      -- CP-element group 57: 	 branch_block_stmt_1642/assign_stmt_1916_to_assign_stmt_1951__entry__
      -- CP-element group 57: 	 branch_block_stmt_1642/if_stmt_1896_else_link/$exit
      -- CP-element group 57: 	 branch_block_stmt_1642/if_stmt_1896_else_link/else_choice_transition
      -- CP-element group 57: 	 branch_block_stmt_1642/whilex_xbody_ifx_xelse
      -- CP-element group 57: 	 branch_block_stmt_1642/assign_stmt_1916_to_assign_stmt_1951/$entry
      -- CP-element group 57: 	 branch_block_stmt_1642/assign_stmt_1916_to_assign_stmt_1951/type_cast_1920_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_1642/assign_stmt_1916_to_assign_stmt_1951/type_cast_1920_update_start_
      -- CP-element group 57: 	 branch_block_stmt_1642/assign_stmt_1916_to_assign_stmt_1951/type_cast_1920_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_1642/assign_stmt_1916_to_assign_stmt_1951/type_cast_1920_Sample/rr
      -- CP-element group 57: 	 branch_block_stmt_1642/assign_stmt_1916_to_assign_stmt_1951/type_cast_1920_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_1642/assign_stmt_1916_to_assign_stmt_1951/type_cast_1920_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_1642/assign_stmt_1916_to_assign_stmt_1951/type_cast_1935_update_start_
      -- CP-element group 57: 	 branch_block_stmt_1642/assign_stmt_1916_to_assign_stmt_1951/type_cast_1935_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_1642/assign_stmt_1916_to_assign_stmt_1951/type_cast_1935_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_1642/assign_stmt_1916_to_assign_stmt_1951/type_cast_1945_update_start_
      -- CP-element group 57: 	 branch_block_stmt_1642/assign_stmt_1916_to_assign_stmt_1951/type_cast_1945_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_1642/assign_stmt_1916_to_assign_stmt_1951/type_cast_1945_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_1642/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 57: 	 branch_block_stmt_1642/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 57: 	 branch_block_stmt_1642/merge_stmt_1910_PhiReqMerge
      -- CP-element group 57: 	 branch_block_stmt_1642/merge_stmt_1910_PhiAck/$entry
      -- CP-element group 57: 	 branch_block_stmt_1642/merge_stmt_1910_PhiAck/$exit
      -- CP-element group 57: 	 branch_block_stmt_1642/merge_stmt_1910_PhiAck/dummy
      -- 
    else_choice_transition_4671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1896_branch_ack_0, ack => convTransposeB_CP_4133_elements(57)); -- 
    rr_4687_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4687_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(57), ack => type_cast_1920_inst_req_0); -- 
    cr_4692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(57), ack => type_cast_1920_inst_req_1); -- 
    cr_4706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(57), ack => type_cast_1935_inst_req_1); -- 
    cr_4720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(57), ack => type_cast_1945_inst_req_1); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_1642/assign_stmt_1916_to_assign_stmt_1951/type_cast_1920_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_1642/assign_stmt_1916_to_assign_stmt_1951/type_cast_1920_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_1642/assign_stmt_1916_to_assign_stmt_1951/type_cast_1920_Sample/ra
      -- 
    ra_4688_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1920_inst_ack_0, ack => convTransposeB_CP_4133_elements(58)); -- 
    -- CP-element group 59:  transition  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (6) 
      -- CP-element group 59: 	 branch_block_stmt_1642/assign_stmt_1916_to_assign_stmt_1951/type_cast_1920_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_1642/assign_stmt_1916_to_assign_stmt_1951/type_cast_1920_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_1642/assign_stmt_1916_to_assign_stmt_1951/type_cast_1920_Update/ca
      -- CP-element group 59: 	 branch_block_stmt_1642/assign_stmt_1916_to_assign_stmt_1951/type_cast_1935_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_1642/assign_stmt_1916_to_assign_stmt_1951/type_cast_1935_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_1642/assign_stmt_1916_to_assign_stmt_1951/type_cast_1935_Sample/rr
      -- 
    ca_4693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1920_inst_ack_1, ack => convTransposeB_CP_4133_elements(59)); -- 
    rr_4701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(59), ack => type_cast_1935_inst_req_0); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_1642/assign_stmt_1916_to_assign_stmt_1951/type_cast_1935_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_1642/assign_stmt_1916_to_assign_stmt_1951/type_cast_1935_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_1642/assign_stmt_1916_to_assign_stmt_1951/type_cast_1935_Sample/ra
      -- 
    ra_4702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1935_inst_ack_0, ack => convTransposeB_CP_4133_elements(60)); -- 
    -- CP-element group 61:  transition  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	57 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_1642/assign_stmt_1916_to_assign_stmt_1951/type_cast_1935_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_1642/assign_stmt_1916_to_assign_stmt_1951/type_cast_1935_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_1642/assign_stmt_1916_to_assign_stmt_1951/type_cast_1935_Update/ca
      -- CP-element group 61: 	 branch_block_stmt_1642/assign_stmt_1916_to_assign_stmt_1951/type_cast_1945_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_1642/assign_stmt_1916_to_assign_stmt_1951/type_cast_1945_Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_1642/assign_stmt_1916_to_assign_stmt_1951/type_cast_1945_Sample/rr
      -- 
    ca_4707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1935_inst_ack_1, ack => convTransposeB_CP_4133_elements(61)); -- 
    rr_4715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(61), ack => type_cast_1945_inst_req_0); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_1642/assign_stmt_1916_to_assign_stmt_1951/type_cast_1945_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_1642/assign_stmt_1916_to_assign_stmt_1951/type_cast_1945_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_1642/assign_stmt_1916_to_assign_stmt_1951/type_cast_1945_Sample/ra
      -- 
    ra_4716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1945_inst_ack_0, ack => convTransposeB_CP_4133_elements(62)); -- 
    -- CP-element group 63:  branch  transition  place  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (13) 
      -- CP-element group 63: 	 branch_block_stmt_1642/assign_stmt_1916_to_assign_stmt_1951__exit__
      -- CP-element group 63: 	 branch_block_stmt_1642/if_stmt_1952__entry__
      -- CP-element group 63: 	 branch_block_stmt_1642/assign_stmt_1916_to_assign_stmt_1951/$exit
      -- CP-element group 63: 	 branch_block_stmt_1642/assign_stmt_1916_to_assign_stmt_1951/type_cast_1945_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_1642/assign_stmt_1916_to_assign_stmt_1951/type_cast_1945_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_1642/assign_stmt_1916_to_assign_stmt_1951/type_cast_1945_Update/ca
      -- CP-element group 63: 	 branch_block_stmt_1642/if_stmt_1952_dead_link/$entry
      -- CP-element group 63: 	 branch_block_stmt_1642/if_stmt_1952_eval_test/$entry
      -- CP-element group 63: 	 branch_block_stmt_1642/if_stmt_1952_eval_test/$exit
      -- CP-element group 63: 	 branch_block_stmt_1642/if_stmt_1952_eval_test/branch_req
      -- CP-element group 63: 	 branch_block_stmt_1642/R_cmp132_1953_place
      -- CP-element group 63: 	 branch_block_stmt_1642/if_stmt_1952_if_link/$entry
      -- CP-element group 63: 	 branch_block_stmt_1642/if_stmt_1952_else_link/$entry
      -- 
    ca_4721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1945_inst_ack_1, ack => convTransposeB_CP_4133_elements(63)); -- 
    branch_req_4729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(63), ack => if_stmt_1952_branch_req_0); -- 
    -- CP-element group 64:  merge  transition  place  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (15) 
      -- CP-element group 64: 	 branch_block_stmt_1642/merge_stmt_1958__exit__
      -- CP-element group 64: 	 branch_block_stmt_1642/assign_stmt_1963__entry__
      -- CP-element group 64: 	 branch_block_stmt_1642/if_stmt_1952_if_link/$exit
      -- CP-element group 64: 	 branch_block_stmt_1642/if_stmt_1952_if_link/if_choice_transition
      -- CP-element group 64: 	 branch_block_stmt_1642/ifx_xelse_whilex_xend
      -- CP-element group 64: 	 branch_block_stmt_1642/assign_stmt_1963/$entry
      -- CP-element group 64: 	 branch_block_stmt_1642/assign_stmt_1963/WPIPE_Block1_done_1960_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_1642/assign_stmt_1963/WPIPE_Block1_done_1960_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_1642/assign_stmt_1963/WPIPE_Block1_done_1960_Sample/req
      -- CP-element group 64: 	 branch_block_stmt_1642/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 64: 	 branch_block_stmt_1642/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 64: 	 branch_block_stmt_1642/merge_stmt_1958_PhiReqMerge
      -- CP-element group 64: 	 branch_block_stmt_1642/merge_stmt_1958_PhiAck/$entry
      -- CP-element group 64: 	 branch_block_stmt_1642/merge_stmt_1958_PhiAck/$exit
      -- CP-element group 64: 	 branch_block_stmt_1642/merge_stmt_1958_PhiAck/dummy
      -- 
    if_choice_transition_4734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1952_branch_ack_1, ack => convTransposeB_CP_4133_elements(64)); -- 
    req_4751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(64), ack => WPIPE_Block1_done_1960_inst_req_0); -- 
    -- CP-element group 65:  fork  transition  place  input  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	73 
    -- CP-element group 65: 	74 
    -- CP-element group 65: 	76 
    -- CP-element group 65: 	77 
    -- CP-element group 65:  members (20) 
      -- CP-element group 65: 	 branch_block_stmt_1642/if_stmt_1952_else_link/$exit
      -- CP-element group 65: 	 branch_block_stmt_1642/if_stmt_1952_else_link/else_choice_transition
      -- CP-element group 65: 	 branch_block_stmt_1642/ifx_xelse_whilex_xbodyx_xouter
      -- CP-element group 65: 	 branch_block_stmt_1642/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 65: 	 branch_block_stmt_1642/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1728/$entry
      -- CP-element group 65: 	 branch_block_stmt_1642/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/$entry
      -- CP-element group 65: 	 branch_block_stmt_1642/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1733/$entry
      -- CP-element group 65: 	 branch_block_stmt_1642/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1733/SplitProtocol/$entry
      -- CP-element group 65: 	 branch_block_stmt_1642/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1733/SplitProtocol/Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_1642/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1733/SplitProtocol/Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_1642/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1733/SplitProtocol/Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1642/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1733/SplitProtocol/Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1642/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/$entry
      -- CP-element group 65: 	 branch_block_stmt_1642/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/$entry
      -- CP-element group 65: 	 branch_block_stmt_1642/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/type_cast_1740/$entry
      -- CP-element group 65: 	 branch_block_stmt_1642/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/type_cast_1740/SplitProtocol/$entry
      -- CP-element group 65: 	 branch_block_stmt_1642/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/type_cast_1740/SplitProtocol/Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_1642/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/type_cast_1740/SplitProtocol/Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_1642/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/type_cast_1740/SplitProtocol/Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1642/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/type_cast_1740/SplitProtocol/Update/cr
      -- 
    else_choice_transition_4738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1952_branch_ack_0, ack => convTransposeB_CP_4133_elements(65)); -- 
    rr_4810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(65), ack => type_cast_1733_inst_req_0); -- 
    cr_4815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(65), ack => type_cast_1733_inst_req_1); -- 
    rr_4833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(65), ack => type_cast_1740_inst_req_0); -- 
    cr_4838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(65), ack => type_cast_1740_inst_req_1); -- 
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_1642/assign_stmt_1963/WPIPE_Block1_done_1960_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_1642/assign_stmt_1963/WPIPE_Block1_done_1960_update_start_
      -- CP-element group 66: 	 branch_block_stmt_1642/assign_stmt_1963/WPIPE_Block1_done_1960_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_1642/assign_stmt_1963/WPIPE_Block1_done_1960_Sample/ack
      -- CP-element group 66: 	 branch_block_stmt_1642/assign_stmt_1963/WPIPE_Block1_done_1960_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_1642/assign_stmt_1963/WPIPE_Block1_done_1960_Update/req
      -- 
    ack_4752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_1960_inst_ack_0, ack => convTransposeB_CP_4133_elements(66)); -- 
    req_4756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(66), ack => WPIPE_Block1_done_1960_inst_req_1); -- 
    -- CP-element group 67:  transition  place  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (16) 
      -- CP-element group 67: 	 branch_block_stmt_1642/merge_stmt_1965__exit__
      -- CP-element group 67: 	 $exit
      -- CP-element group 67: 	 branch_block_stmt_1642/$exit
      -- CP-element group 67: 	 branch_block_stmt_1642/branch_block_stmt_1642__exit__
      -- CP-element group 67: 	 branch_block_stmt_1642/assign_stmt_1963__exit__
      -- CP-element group 67: 	 branch_block_stmt_1642/return__
      -- CP-element group 67: 	 branch_block_stmt_1642/assign_stmt_1963/$exit
      -- CP-element group 67: 	 branch_block_stmt_1642/assign_stmt_1963/WPIPE_Block1_done_1960_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_1642/assign_stmt_1963/WPIPE_Block1_done_1960_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_1642/assign_stmt_1963/WPIPE_Block1_done_1960_Update/ack
      -- CP-element group 67: 	 branch_block_stmt_1642/return___PhiReq/$entry
      -- CP-element group 67: 	 branch_block_stmt_1642/return___PhiReq/$exit
      -- CP-element group 67: 	 branch_block_stmt_1642/merge_stmt_1965_PhiReqMerge
      -- CP-element group 67: 	 branch_block_stmt_1642/merge_stmt_1965_PhiAck/$entry
      -- CP-element group 67: 	 branch_block_stmt_1642/merge_stmt_1965_PhiAck/$exit
      -- CP-element group 67: 	 branch_block_stmt_1642/merge_stmt_1965_PhiAck/dummy
      -- 
    ack_4757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_1960_inst_ack_1, ack => convTransposeB_CP_4133_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	31 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (2) 
      -- CP-element group 68: 	 branch_block_stmt_1642/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1731/SplitProtocol/Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_1642/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1731/SplitProtocol/Sample/ra
      -- 
    ra_4777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1731_inst_ack_0, ack => convTransposeB_CP_4133_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	31 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (2) 
      -- CP-element group 69: 	 branch_block_stmt_1642/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1731/SplitProtocol/Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_1642/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1731/SplitProtocol/Update/ca
      -- 
    ca_4782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1731_inst_ack_1, ack => convTransposeB_CP_4133_elements(69)); -- 
    -- CP-element group 70:  join  transition  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (5) 
      -- CP-element group 70: 	 branch_block_stmt_1642/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1728/$exit
      -- CP-element group 70: 	 branch_block_stmt_1642/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/$exit
      -- CP-element group 70: 	 branch_block_stmt_1642/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1731/$exit
      -- CP-element group 70: 	 branch_block_stmt_1642/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1731/SplitProtocol/$exit
      -- CP-element group 70: 	 branch_block_stmt_1642/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1728/phi_stmt_1728_req
      -- 
    phi_stmt_1728_req_4783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1728_req_4783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(70), ack => phi_stmt_1728_req_0); -- 
    convTransposeB_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4133_elements(68) & convTransposeB_CP_4133_elements(69);
      gj_convTransposeB_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4133_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  transition  output  delay-element  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	31 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (4) 
      -- CP-element group 71: 	 branch_block_stmt_1642/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/$exit
      -- CP-element group 71: 	 branch_block_stmt_1642/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/$exit
      -- CP-element group 71: 	 branch_block_stmt_1642/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/type_cast_1738_konst_delay_trans
      -- CP-element group 71: 	 branch_block_stmt_1642/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_req
      -- 
    phi_stmt_1734_req_4791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1734_req_4791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(71), ack => phi_stmt_1734_req_0); -- 
    -- Element group convTransposeB_CP_4133_elements(71) is a control-delay.
    cp_element_71_delay: control_delay_element  generic map(name => " 71_delay", delay_value => 1)  port map(req => convTransposeB_CP_4133_elements(31), ack => convTransposeB_CP_4133_elements(71), clk => clk, reset =>reset);
    -- CP-element group 72:  join  transition  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	80 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_1642/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4133_elements(70) & convTransposeB_CP_4133_elements(71);
      gj_convTransposeB_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4133_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	65 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (2) 
      -- CP-element group 73: 	 branch_block_stmt_1642/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1733/SplitProtocol/Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_1642/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1733/SplitProtocol/Sample/ra
      -- 
    ra_4811_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1733_inst_ack_0, ack => convTransposeB_CP_4133_elements(73)); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	65 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74:  members (2) 
      -- CP-element group 74: 	 branch_block_stmt_1642/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1733/SplitProtocol/Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_1642/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1733/SplitProtocol/Update/ca
      -- 
    ca_4816_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1733_inst_ack_1, ack => convTransposeB_CP_4133_elements(74)); -- 
    -- CP-element group 75:  join  transition  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	79 
    -- CP-element group 75:  members (5) 
      -- CP-element group 75: 	 branch_block_stmt_1642/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1728/$exit
      -- CP-element group 75: 	 branch_block_stmt_1642/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/$exit
      -- CP-element group 75: 	 branch_block_stmt_1642/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1733/$exit
      -- CP-element group 75: 	 branch_block_stmt_1642/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1733/SplitProtocol/$exit
      -- CP-element group 75: 	 branch_block_stmt_1642/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1728/phi_stmt_1728_req
      -- 
    phi_stmt_1728_req_4817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1728_req_4817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(75), ack => phi_stmt_1728_req_1); -- 
    convTransposeB_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4133_elements(73) & convTransposeB_CP_4133_elements(74);
      gj_convTransposeB_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4133_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	65 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (2) 
      -- CP-element group 76: 	 branch_block_stmt_1642/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/type_cast_1740/SplitProtocol/Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_1642/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/type_cast_1740/SplitProtocol/Sample/ra
      -- 
    ra_4834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1740_inst_ack_0, ack => convTransposeB_CP_4133_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	65 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_1642/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/type_cast_1740/SplitProtocol/Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_1642/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/type_cast_1740/SplitProtocol/Update/ca
      -- 
    ca_4839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1740_inst_ack_1, ack => convTransposeB_CP_4133_elements(77)); -- 
    -- CP-element group 78:  join  transition  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (5) 
      -- CP-element group 78: 	 branch_block_stmt_1642/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/$exit
      -- CP-element group 78: 	 branch_block_stmt_1642/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/$exit
      -- CP-element group 78: 	 branch_block_stmt_1642/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/type_cast_1740/$exit
      -- CP-element group 78: 	 branch_block_stmt_1642/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/type_cast_1740/SplitProtocol/$exit
      -- CP-element group 78: 	 branch_block_stmt_1642/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_req
      -- 
    phi_stmt_1734_req_4840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1734_req_4840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(78), ack => phi_stmt_1734_req_1); -- 
    convTransposeB_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4133_elements(76) & convTransposeB_CP_4133_elements(77);
      gj_convTransposeB_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4133_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  join  transition  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	75 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_1642/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4133_elements(75) & convTransposeB_CP_4133_elements(78);
      gj_convTransposeB_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4133_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  merge  fork  transition  place  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	72 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_1642/merge_stmt_1727_PhiReqMerge
      -- CP-element group 80: 	 branch_block_stmt_1642/merge_stmt_1727_PhiAck/$entry
      -- 
    convTransposeB_CP_4133_elements(80) <= OrReduce(convTransposeB_CP_4133_elements(72) & convTransposeB_CP_4133_elements(79));
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_1642/merge_stmt_1727_PhiAck/phi_stmt_1728_ack
      -- 
    phi_stmt_1728_ack_4845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1728_ack_0, ack => convTransposeB_CP_4133_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_1642/merge_stmt_1727_PhiAck/phi_stmt_1734_ack
      -- 
    phi_stmt_1734_ack_4846_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1734_ack_0, ack => convTransposeB_CP_4133_elements(82)); -- 
    -- CP-element group 83:  join  transition  place  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	87 
    -- CP-element group 83:  members (10) 
      -- CP-element group 83: 	 branch_block_stmt_1642/assign_stmt_1746_to_assign_stmt_1791/$entry
      -- CP-element group 83: 	 branch_block_stmt_1642/assign_stmt_1746_to_assign_stmt_1791/$exit
      -- CP-element group 83: 	 branch_block_stmt_1642/merge_stmt_1727__exit__
      -- CP-element group 83: 	 branch_block_stmt_1642/assign_stmt_1746_to_assign_stmt_1791__entry__
      -- CP-element group 83: 	 branch_block_stmt_1642/assign_stmt_1746_to_assign_stmt_1791__exit__
      -- CP-element group 83: 	 branch_block_stmt_1642/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 83: 	 branch_block_stmt_1642/merge_stmt_1727_PhiAck/$exit
      -- CP-element group 83: 	 branch_block_stmt_1642/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- CP-element group 83: 	 branch_block_stmt_1642/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1794/$entry
      -- CP-element group 83: 	 branch_block_stmt_1642/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/$entry
      -- 
    convTransposeB_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4133_elements(81) & convTransposeB_CP_4133_elements(82);
      gj_convTransposeB_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4133_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	56 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_1642/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/type_cast_1797/SplitProtocol/Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_1642/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/type_cast_1797/SplitProtocol/Sample/ra
      -- 
    ra_4866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1797_inst_ack_0, ack => convTransposeB_CP_4133_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	56 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_1642/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/type_cast_1797/SplitProtocol/Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_1642/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/type_cast_1797/SplitProtocol/Update/ca
      -- 
    ca_4871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1797_inst_ack_1, ack => convTransposeB_CP_4133_elements(85)); -- 
    -- CP-element group 86:  join  transition  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (6) 
      -- CP-element group 86: 	 branch_block_stmt_1642/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- CP-element group 86: 	 branch_block_stmt_1642/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1794/$exit
      -- CP-element group 86: 	 branch_block_stmt_1642/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/$exit
      -- CP-element group 86: 	 branch_block_stmt_1642/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/type_cast_1797/$exit
      -- CP-element group 86: 	 branch_block_stmt_1642/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/type_cast_1797/SplitProtocol/$exit
      -- CP-element group 86: 	 branch_block_stmt_1642/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1794/phi_stmt_1794_req
      -- 
    phi_stmt_1794_req_4872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1794_req_4872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(86), ack => phi_stmt_1794_req_0); -- 
    convTransposeB_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4133_elements(84) & convTransposeB_CP_4133_elements(85);
      gj_convTransposeB_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4133_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  transition  output  delay-element  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	83 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (5) 
      -- CP-element group 87: 	 branch_block_stmt_1642/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- CP-element group 87: 	 branch_block_stmt_1642/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1794/$exit
      -- CP-element group 87: 	 branch_block_stmt_1642/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/$exit
      -- CP-element group 87: 	 branch_block_stmt_1642/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/type_cast_1800_konst_delay_trans
      -- CP-element group 87: 	 branch_block_stmt_1642/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1794/phi_stmt_1794_req
      -- 
    phi_stmt_1794_req_4883_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1794_req_4883_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(87), ack => phi_stmt_1794_req_1); -- 
    -- Element group convTransposeB_CP_4133_elements(87) is a control-delay.
    cp_element_87_delay: control_delay_element  generic map(name => " 87_delay", delay_value => 1)  port map(req => convTransposeB_CP_4133_elements(83), ack => convTransposeB_CP_4133_elements(87), clk => clk, reset =>reset);
    -- CP-element group 88:  merge  transition  place  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_1642/merge_stmt_1793_PhiReqMerge
      -- CP-element group 88: 	 branch_block_stmt_1642/merge_stmt_1793_PhiAck/$entry
      -- 
    convTransposeB_CP_4133_elements(88) <= OrReduce(convTransposeB_CP_4133_elements(86) & convTransposeB_CP_4133_elements(87));
    -- CP-element group 89:  fork  transition  place  input  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	32 
    -- CP-element group 89: 	33 
    -- CP-element group 89: 	35 
    -- CP-element group 89: 	37 
    -- CP-element group 89: 	39 
    -- CP-element group 89: 	41 
    -- CP-element group 89: 	42 
    -- CP-element group 89: 	43 
    -- CP-element group 89: 	45 
    -- CP-element group 89: 	47 
    -- CP-element group 89: 	49 
    -- CP-element group 89: 	52 
    -- CP-element group 89: 	53 
    -- CP-element group 89: 	54 
    -- CP-element group 89:  members (51) 
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1835_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/$entry
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1821_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1821_Sample/rr
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1821_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1821_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/addr_of_1842_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1835_Update/cr
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1821_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1835_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1821_Update/cr
      -- CP-element group 89: 	 branch_block_stmt_1642/merge_stmt_1793__exit__
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895__entry__
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1841_final_index_sum_regn_update_start
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1841_final_index_sum_regn_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1841_final_index_sum_regn_Update/req
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/addr_of_1842_complete/$entry
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/addr_of_1842_complete/req
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1846_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1846_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1846_Update/word_access_complete/$entry
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1846_Update/word_access_complete/word_0/$entry
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1846_Update/word_access_complete/word_0/cr
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1851_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1851_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1851_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1851_Sample/rr
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1851_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1851_Update/cr
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1865_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1865_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1865_Update/cr
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/addr_of_1872_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1871_final_index_sum_regn_update_start
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1871_final_index_sum_regn_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/array_obj_ref_1871_final_index_sum_regn_Update/req
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/addr_of_1872_complete/$entry
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/addr_of_1872_complete/req
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1875_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1875_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1875_Update/word_access_complete/$entry
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1875_Update/word_access_complete/word_0/$entry
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/ptr_deref_1875_Update/word_access_complete/word_0/cr
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1881_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1881_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1881_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1881_Sample/rr
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1881_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1642/assign_stmt_1807_to_assign_stmt_1895/type_cast_1881_Update/cr
      -- CP-element group 89: 	 branch_block_stmt_1642/merge_stmt_1793_PhiAck/$exit
      -- CP-element group 89: 	 branch_block_stmt_1642/merge_stmt_1793_PhiAck/phi_stmt_1794_ack
      -- 
    phi_stmt_1794_ack_4888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1794_ack_0, ack => convTransposeB_CP_4133_elements(89)); -- 
    rr_4400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(89), ack => type_cast_1821_inst_req_0); -- 
    cr_4419_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4419_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(89), ack => type_cast_1835_inst_req_1); -- 
    cr_4405_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4405_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(89), ack => type_cast_1821_inst_req_1); -- 
    req_4450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(89), ack => array_obj_ref_1841_index_offset_req_1); -- 
    req_4465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(89), ack => addr_of_1842_final_reg_req_1); -- 
    cr_4510_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4510_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(89), ack => ptr_deref_1846_load_0_req_1); -- 
    rr_4524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(89), ack => type_cast_1851_inst_req_0); -- 
    cr_4529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(89), ack => type_cast_1851_inst_req_1); -- 
    cr_4543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(89), ack => type_cast_1865_inst_req_1); -- 
    req_4574_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4574_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(89), ack => array_obj_ref_1871_index_offset_req_1); -- 
    req_4589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(89), ack => addr_of_1872_final_reg_req_1); -- 
    cr_4639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(89), ack => ptr_deref_1875_store_0_req_1); -- 
    rr_4648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(89), ack => type_cast_1881_inst_req_0); -- 
    cr_4653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4133_elements(89), ack => type_cast_1881_inst_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_1829_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1859_wire : std_logic_vector(31 downto 0);
    signal R_idxprom96_1870_resized : std_logic_vector(13 downto 0);
    signal R_idxprom96_1870_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_1840_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_1840_scaled : std_logic_vector(13 downto 0);
    signal add101_1888 : std_logic_vector(31 downto 0);
    signal add43_1812 : std_logic_vector(15 downto 0);
    signal add87_1817 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1841_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1841_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1841_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1841_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1841_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1841_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1871_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1871_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1871_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1871_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1871_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1871_root_address : std_logic_vector(13 downto 0);
    signal arrayidx91_1843 : std_logic_vector(31 downto 0);
    signal arrayidx97_1873 : std_logic_vector(31 downto 0);
    signal call11_1663 : std_logic_vector(15 downto 0);
    signal call13_1666 : std_logic_vector(15 downto 0);
    signal call14_1669 : std_logic_vector(15 downto 0);
    signal call15_1672 : std_logic_vector(15 downto 0);
    signal call17_1675 : std_logic_vector(15 downto 0);
    signal call19_1678 : std_logic_vector(15 downto 0);
    signal call1_1648 : std_logic_vector(15 downto 0);
    signal call3_1651 : std_logic_vector(15 downto 0);
    signal call5_1654 : std_logic_vector(15 downto 0);
    signal call7_1657 : std_logic_vector(15 downto 0);
    signal call9_1660 : std_logic_vector(15 downto 0);
    signal call_1645 : std_logic_vector(15 downto 0);
    signal cmp116_1926 : std_logic_vector(0 downto 0);
    signal cmp132_1951 : std_logic_vector(0 downto 0);
    signal cmp_1895 : std_logic_vector(0 downto 0);
    signal conv100_1882 : std_logic_vector(31 downto 0);
    signal conv104_1689 : std_logic_vector(31 downto 0);
    signal conv112_1921 : std_logic_vector(31 downto 0);
    signal conv115_1693 : std_logic_vector(31 downto 0);
    signal conv127_1946 : std_logic_vector(31 downto 0);
    signal conv130_1697 : std_logic_vector(31 downto 0);
    signal conv90_1822 : std_logic_vector(31 downto 0);
    signal conv94_1852 : std_logic_vector(31 downto 0);
    signal div131_1703 : std_logic_vector(31 downto 0);
    signal div_1685 : std_logic_vector(15 downto 0);
    signal idxprom96_1866 : std_logic_vector(63 downto 0);
    signal idxprom_1836 : std_logic_vector(63 downto 0);
    signal inc120_1936 : std_logic_vector(15 downto 0);
    signal inc_1916 : std_logic_vector(15 downto 0);
    signal indvar_1794 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_1908 : std_logic_vector(15 downto 0);
    signal input_dim0x_x0_1941 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_1734 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_1728 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_1932 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1807 : std_logic_vector(15 downto 0);
    signal ptr_deref_1846_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1846_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1846_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1846_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1846_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1875_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1875_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1875_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1875_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1875_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1875_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr95_1861 : std_logic_vector(31 downto 0);
    signal shr_1831 : std_logic_vector(31 downto 0);
    signal tmp10_1791 : std_logic_vector(15 downto 0);
    signal tmp159_1746 : std_logic_vector(15 downto 0);
    signal tmp160_1751 : std_logic_vector(15 downto 0);
    signal tmp161_1756 : std_logic_vector(15 downto 0);
    signal tmp1_1714 : std_logic_vector(15 downto 0);
    signal tmp2_1761 : std_logic_vector(15 downto 0);
    signal tmp3_1766 : std_logic_vector(15 downto 0);
    signal tmp4_1720 : std_logic_vector(15 downto 0);
    signal tmp5_1725 : std_logic_vector(15 downto 0);
    signal tmp6_1771 : std_logic_vector(15 downto 0);
    signal tmp7_1776 : std_logic_vector(15 downto 0);
    signal tmp8_1781 : std_logic_vector(15 downto 0);
    signal tmp92_1847 : std_logic_vector(63 downto 0);
    signal tmp9_1786 : std_logic_vector(15 downto 0);
    signal tmp_1709 : std_logic_vector(15 downto 0);
    signal type_cast_1683_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1701_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1707_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1718_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1731_wire : std_logic_vector(15 downto 0);
    signal type_cast_1733_wire : std_logic_vector(15 downto 0);
    signal type_cast_1738_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1740_wire : std_logic_vector(15 downto 0);
    signal type_cast_1797_wire : std_logic_vector(15 downto 0);
    signal type_cast_1800_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1805_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1820_wire : std_logic_vector(31 downto 0);
    signal type_cast_1825_wire : std_logic_vector(31 downto 0);
    signal type_cast_1828_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1834_wire : std_logic_vector(63 downto 0);
    signal type_cast_1850_wire : std_logic_vector(31 downto 0);
    signal type_cast_1855_wire : std_logic_vector(31 downto 0);
    signal type_cast_1858_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1864_wire : std_logic_vector(63 downto 0);
    signal type_cast_1880_wire : std_logic_vector(31 downto 0);
    signal type_cast_1886_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1891_wire : std_logic_vector(31 downto 0);
    signal type_cast_1893_wire : std_logic_vector(31 downto 0);
    signal type_cast_1906_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1914_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1919_wire : std_logic_vector(31 downto 0);
    signal type_cast_1944_wire : std_logic_vector(31 downto 0);
    signal type_cast_1962_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_1841_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1841_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1841_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1841_resized_base_address <= "00000000000000";
    array_obj_ref_1871_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1871_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1871_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1871_resized_base_address <= "00000000000000";
    ptr_deref_1846_word_offset_0 <= "00000000000000";
    ptr_deref_1875_word_offset_0 <= "00000000000000";
    type_cast_1683_wire_constant <= "0000000000000001";
    type_cast_1701_wire_constant <= "00000000000000000000000000000001";
    type_cast_1707_wire_constant <= "1111111111111111";
    type_cast_1718_wire_constant <= "1111111111111111";
    type_cast_1738_wire_constant <= "0000000000000000";
    type_cast_1800_wire_constant <= "0000000000000000";
    type_cast_1805_wire_constant <= "0000000000000100";
    type_cast_1828_wire_constant <= "00000000000000000000000000000010";
    type_cast_1858_wire_constant <= "00000000000000000000000000000010";
    type_cast_1886_wire_constant <= "00000000000000000000000000000100";
    type_cast_1906_wire_constant <= "0000000000000001";
    type_cast_1914_wire_constant <= "0000000000000001";
    type_cast_1962_wire_constant <= "0000000000000001";
    phi_stmt_1728: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1731_wire & type_cast_1733_wire;
      req <= phi_stmt_1728_req_0 & phi_stmt_1728_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1728",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1728_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_1728,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1728
    phi_stmt_1734: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1738_wire_constant & type_cast_1740_wire;
      req <= phi_stmt_1734_req_0 & phi_stmt_1734_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1734",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1734_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_1734,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1734
    phi_stmt_1794: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1797_wire & type_cast_1800_wire_constant;
      req <= phi_stmt_1794_req_0 & phi_stmt_1794_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1794",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1794_ack_0,
          idata => idata,
          odata => indvar_1794,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1794
    -- flow-through select operator MUX_1931_inst
    input_dim1x_x2_1932 <= div_1685 when (cmp116_1926(0) /=  '0') else inc_1916;
    addr_of_1842_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1842_final_reg_req_0;
      addr_of_1842_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1842_final_reg_req_1;
      addr_of_1842_final_reg_ack_1<= rack(0);
      addr_of_1842_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1842_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1841_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx91_1843,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1872_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1872_final_reg_req_0;
      addr_of_1872_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1872_final_reg_req_1;
      addr_of_1872_final_reg_ack_1<= rack(0);
      addr_of_1872_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1872_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1871_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx97_1873,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1688_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1688_inst_req_0;
      type_cast_1688_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1688_inst_req_1;
      type_cast_1688_inst_ack_1<= rack(0);
      type_cast_1688_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1688_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_1651,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv104_1689,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1692_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1692_inst_req_0;
      type_cast_1692_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1692_inst_req_1;
      type_cast_1692_inst_ack_1<= rack(0);
      type_cast_1692_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1692_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1_1648,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv115_1693,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1696_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1696_inst_req_0;
      type_cast_1696_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1696_inst_req_1;
      type_cast_1696_inst_ack_1<= rack(0);
      type_cast_1696_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1696_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1645,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv130_1697,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1731_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1731_inst_req_0;
      type_cast_1731_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1731_inst_req_1;
      type_cast_1731_inst_ack_1<= rack(0);
      type_cast_1731_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1731_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_1685,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1731_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1733_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1733_inst_req_0;
      type_cast_1733_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1733_inst_req_1;
      type_cast_1733_inst_ack_1<= rack(0);
      type_cast_1733_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1733_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_1932,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1733_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1740_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1740_inst_req_0;
      type_cast_1740_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1740_inst_req_1;
      type_cast_1740_inst_ack_1<= rack(0);
      type_cast_1740_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1740_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x0_1941,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1740_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1797_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1797_inst_req_0;
      type_cast_1797_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1797_inst_req_1;
      type_cast_1797_inst_ack_1<= rack(0);
      type_cast_1797_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1797_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1908,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1797_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1821_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1821_inst_req_0;
      type_cast_1821_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1821_inst_req_1;
      type_cast_1821_inst_ack_1<= rack(0);
      type_cast_1821_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1821_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1820_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_1822,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1825_inst
    process(conv90_1822) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv90_1822(31 downto 0);
      type_cast_1825_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1830_inst
    process(ASHR_i32_i32_1829_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1829_wire(31 downto 0);
      shr_1831 <= tmp_var; -- 
    end process;
    type_cast_1835_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1835_inst_req_0;
      type_cast_1835_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1835_inst_req_1;
      type_cast_1835_inst_ack_1<= rack(0);
      type_cast_1835_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1835_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1834_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_1836,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1851_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1851_inst_req_0;
      type_cast_1851_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1851_inst_req_1;
      type_cast_1851_inst_ack_1<= rack(0);
      type_cast_1851_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1851_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1850_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv94_1852,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1855_inst
    process(conv94_1852) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv94_1852(31 downto 0);
      type_cast_1855_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1860_inst
    process(ASHR_i32_i32_1859_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1859_wire(31 downto 0);
      shr95_1861 <= tmp_var; -- 
    end process;
    type_cast_1865_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1865_inst_req_0;
      type_cast_1865_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1865_inst_req_1;
      type_cast_1865_inst_ack_1<= rack(0);
      type_cast_1865_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1865_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1864_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom96_1866,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1881_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1881_inst_req_0;
      type_cast_1881_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1881_inst_req_1;
      type_cast_1881_inst_ack_1<= rack(0);
      type_cast_1881_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1881_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1880_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv100_1882,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1891_inst
    process(add101_1888) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add101_1888(31 downto 0);
      type_cast_1891_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1893_inst
    process(conv104_1689) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv104_1689(31 downto 0);
      type_cast_1893_wire <= tmp_var; -- 
    end process;
    type_cast_1920_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1920_inst_req_0;
      type_cast_1920_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1920_inst_req_1;
      type_cast_1920_inst_ack_1<= rack(0);
      type_cast_1920_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1920_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1919_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv112_1921,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1935_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1935_inst_req_0;
      type_cast_1935_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1935_inst_req_1;
      type_cast_1935_inst_ack_1<= rack(0);
      type_cast_1935_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1935_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp116_1926,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc120_1936,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1945_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1945_inst_req_0;
      type_cast_1945_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1945_inst_req_1;
      type_cast_1945_inst_ack_1<= rack(0);
      type_cast_1945_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1945_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1944_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv127_1946,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1841_index_1_rename
    process(R_idxprom_1840_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_1840_resized;
      ov(13 downto 0) := iv;
      R_idxprom_1840_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1841_index_1_resize
    process(idxprom_1836) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_1836;
      ov := iv(13 downto 0);
      R_idxprom_1840_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1841_root_address_inst
    process(array_obj_ref_1841_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1841_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1841_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1871_index_1_rename
    process(R_idxprom96_1870_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom96_1870_resized;
      ov(13 downto 0) := iv;
      R_idxprom96_1870_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1871_index_1_resize
    process(idxprom96_1866) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom96_1866;
      ov := iv(13 downto 0);
      R_idxprom96_1870_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1871_root_address_inst
    process(array_obj_ref_1871_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1871_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1871_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1846_addr_0
    process(ptr_deref_1846_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1846_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1846_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1846_base_resize
    process(arrayidx91_1843) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx91_1843;
      ov := iv(13 downto 0);
      ptr_deref_1846_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1846_gather_scatter
    process(ptr_deref_1846_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1846_data_0;
      ov(63 downto 0) := iv;
      tmp92_1847 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1846_root_address_inst
    process(ptr_deref_1846_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1846_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1846_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1875_addr_0
    process(ptr_deref_1875_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1875_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1875_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1875_base_resize
    process(arrayidx97_1873) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx97_1873;
      ov := iv(13 downto 0);
      ptr_deref_1875_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1875_gather_scatter
    process(tmp92_1847) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp92_1847;
      ov(63 downto 0) := iv;
      ptr_deref_1875_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1875_root_address_inst
    process(ptr_deref_1875_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1875_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1875_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1896_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_1895;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1896_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1896_branch_req_0,
          ack0 => if_stmt_1896_branch_ack_0,
          ack1 => if_stmt_1896_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1952_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp132_1951;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1952_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1952_branch_req_0,
          ack0 => if_stmt_1952_branch_ack_0,
          ack1 => if_stmt_1952_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1708_inst
    process(call9_1660) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_1660, type_cast_1707_wire_constant, tmp_var);
      tmp_1709 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1719_inst
    process(call7_1657) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_1657, type_cast_1718_wire_constant, tmp_var);
      tmp4_1720 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1750_inst
    process(input_dim1x_x1x_xph_1728, tmp159_1746) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_1728, tmp159_1746, tmp_var);
      tmp160_1751 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1765_inst
    process(tmp1_1714, tmp2_1761) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp1_1714, tmp2_1761, tmp_var);
      tmp3_1766 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1775_inst
    process(tmp5_1725, tmp6_1771) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp5_1725, tmp6_1771, tmp_var);
      tmp7_1776 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1785_inst
    process(tmp3_1766, tmp8_1781) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp3_1766, tmp8_1781, tmp_var);
      tmp9_1786 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1811_inst
    process(tmp161_1756, input_dim2x_x1_1807) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp161_1756, input_dim2x_x1_1807, tmp_var);
      add43_1812 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1816_inst
    process(tmp10_1791, input_dim2x_x1_1807) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp10_1791, input_dim2x_x1_1807, tmp_var);
      add87_1817 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1907_inst
    process(indvar_1794) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1794, type_cast_1906_wire_constant, tmp_var);
      indvarx_xnext_1908 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1915_inst
    process(input_dim1x_x1x_xph_1728) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_1728, type_cast_1914_wire_constant, tmp_var);
      inc_1916 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1940_inst
    process(inc120_1936, input_dim0x_x2x_xph_1734) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc120_1936, input_dim0x_x2x_xph_1734, tmp_var);
      input_dim0x_x0_1941 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1887_inst
    process(conv100_1882) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv100_1882, type_cast_1886_wire_constant, tmp_var);
      add101_1888 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1829_inst
    process(type_cast_1825_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1825_wire, type_cast_1828_wire_constant, tmp_var);
      ASHR_i32_i32_1829_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1859_inst
    process(type_cast_1855_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1855_wire, type_cast_1858_wire_constant, tmp_var);
      ASHR_i32_i32_1859_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1925_inst
    process(conv112_1921, conv115_1693) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv112_1921, conv115_1693, tmp_var);
      cmp116_1926 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1950_inst
    process(conv127_1946, div131_1703) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv127_1946, div131_1703, tmp_var);
      cmp132_1951 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_1684_inst
    process(call1_1648) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call1_1648, type_cast_1683_wire_constant, tmp_var);
      div_1685 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1702_inst
    process(conv130_1697) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv130_1697, type_cast_1701_wire_constant, tmp_var);
      div131_1703 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1745_inst
    process(call1_1648, input_dim0x_x2x_xph_1734) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call1_1648, input_dim0x_x2x_xph_1734, tmp_var);
      tmp159_1746 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1755_inst
    process(call3_1651, tmp160_1751) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call3_1651, tmp160_1751, tmp_var);
      tmp161_1756 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1760_inst
    process(call13_1666, input_dim1x_x1x_xph_1728) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call13_1666, input_dim1x_x1x_xph_1728, tmp_var);
      tmp2_1761 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1770_inst
    process(call13_1666, input_dim0x_x2x_xph_1734) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call13_1666, input_dim0x_x2x_xph_1734, tmp_var);
      tmp6_1771 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1780_inst
    process(call17_1675, tmp7_1776) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call17_1675, tmp7_1776, tmp_var);
      tmp8_1781 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1790_inst
    process(call19_1678, tmp9_1786) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call19_1678, tmp9_1786, tmp_var);
      tmp10_1791 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1806_inst
    process(indvar_1794) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_1794, type_cast_1805_wire_constant, tmp_var);
      input_dim2x_x1_1807 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1894_inst
    process(type_cast_1891_wire, type_cast_1893_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1891_wire, type_cast_1893_wire, tmp_var);
      cmp_1895 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1713_inst
    process(tmp_1709, call14_1669) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp_1709, call14_1669, tmp_var);
      tmp1_1714 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1724_inst
    process(tmp4_1720, call14_1669) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp4_1720, call14_1669, tmp_var);
      tmp5_1725 <= tmp_var; --
    end process;
    -- shared split operator group (28) : array_obj_ref_1841_index_offset 
    ApIntAdd_group_28: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_1840_scaled;
      array_obj_ref_1841_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1841_index_offset_req_0;
      array_obj_ref_1841_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1841_index_offset_req_1;
      array_obj_ref_1841_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_28_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_28_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : array_obj_ref_1871_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom96_1870_scaled;
      array_obj_ref_1871_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1871_index_offset_req_0;
      array_obj_ref_1871_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1871_index_offset_req_1;
      array_obj_ref_1871_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- unary operator type_cast_1820_inst
    process(add43_1812) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", add43_1812, tmp_var);
      type_cast_1820_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1834_inst
    process(shr_1831) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_1831, tmp_var);
      type_cast_1834_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1850_inst
    process(add87_1817) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", add87_1817, tmp_var);
      type_cast_1850_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1864_inst
    process(shr95_1861) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr95_1861, tmp_var);
      type_cast_1864_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1880_inst
    process(input_dim2x_x1_1807) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim2x_x1_1807, tmp_var);
      type_cast_1880_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1919_inst
    process(inc_1916) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_1916, tmp_var);
      type_cast_1919_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1944_inst
    process(input_dim0x_x0_1941) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim0x_x0_1941, tmp_var);
      type_cast_1944_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_1846_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1846_load_0_req_0;
      ptr_deref_1846_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1846_load_0_req_1;
      ptr_deref_1846_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1846_word_address_0;
      ptr_deref_1846_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_1875_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1875_store_0_req_0;
      ptr_deref_1875_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1875_store_0_req_1;
      ptr_deref_1875_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1875_word_address_0;
      data_in <= ptr_deref_1875_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block1_start_1644_inst RPIPE_Block1_start_1647_inst RPIPE_Block1_start_1650_inst RPIPE_Block1_start_1653_inst RPIPE_Block1_start_1656_inst RPIPE_Block1_start_1659_inst RPIPE_Block1_start_1662_inst RPIPE_Block1_start_1665_inst RPIPE_Block1_start_1668_inst RPIPE_Block1_start_1671_inst RPIPE_Block1_start_1674_inst RPIPE_Block1_start_1677_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(191 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 11 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 11 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 11 downto 0);
      signal guard_vector : std_logic_vector( 11 downto 0);
      constant outBUFs : IntegerArray(11 downto 0) := (11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(11 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false);
      constant guardBuffering: IntegerArray(11 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2);
      -- 
    begin -- 
      reqL_unguarded(11) <= RPIPE_Block1_start_1644_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block1_start_1647_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block1_start_1650_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block1_start_1653_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block1_start_1656_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block1_start_1659_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block1_start_1662_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block1_start_1665_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block1_start_1668_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block1_start_1671_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block1_start_1674_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block1_start_1677_inst_req_0;
      RPIPE_Block1_start_1644_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block1_start_1647_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block1_start_1650_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block1_start_1653_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block1_start_1656_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block1_start_1659_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block1_start_1662_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block1_start_1665_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block1_start_1668_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block1_start_1671_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block1_start_1674_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block1_start_1677_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(11) <= RPIPE_Block1_start_1644_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block1_start_1647_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block1_start_1650_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block1_start_1653_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block1_start_1656_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block1_start_1659_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block1_start_1662_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block1_start_1665_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block1_start_1668_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block1_start_1671_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block1_start_1674_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block1_start_1677_inst_req_1;
      RPIPE_Block1_start_1644_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block1_start_1647_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block1_start_1650_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block1_start_1653_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block1_start_1656_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block1_start_1659_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block1_start_1662_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block1_start_1665_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block1_start_1668_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block1_start_1671_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block1_start_1674_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block1_start_1677_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      call_1645 <= data_out(191 downto 176);
      call1_1648 <= data_out(175 downto 160);
      call3_1651 <= data_out(159 downto 144);
      call5_1654 <= data_out(143 downto 128);
      call7_1657 <= data_out(127 downto 112);
      call9_1660 <= data_out(111 downto 96);
      call11_1663 <= data_out(95 downto 80);
      call13_1666 <= data_out(79 downto 64);
      call14_1669 <= data_out(63 downto 48);
      call15_1672 <= data_out(47 downto 32);
      call17_1675 <= data_out(31 downto 16);
      call19_1678 <= data_out(15 downto 0);
      Block1_start_read_0_gI: SplitGuardInterface generic map(name => "Block1_start_read_0_gI", nreqs => 12, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_start_read_0: InputPortRevised -- 
        generic map ( name => "Block1_start_read_0", data_width => 16,  num_reqs => 12,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_start_pipe_read_req(0),
          oack => Block1_start_pipe_read_ack(0),
          odata => Block1_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block1_done_1960_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block1_done_1960_inst_req_0;
      WPIPE_Block1_done_1960_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block1_done_1960_inst_req_1;
      WPIPE_Block1_done_1960_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_1962_wire_constant;
      Block1_done_write_0_gI: SplitGuardInterface generic map(name => "Block1_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block1_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_done_pipe_write_req(0),
          oack => Block1_done_pipe_write_ack(0),
          odata => Block1_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeB_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeC is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeC;
architecture convTransposeC_arch of convTransposeC is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeC_CP_4929_start: Boolean;
  signal convTransposeC_CP_4929_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal array_obj_ref_2168_index_offset_ack_0 : boolean;
  signal array_obj_ref_2168_index_offset_req_1 : boolean;
  signal type_cast_2178_inst_req_1 : boolean;
  signal type_cast_2065_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1971_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1971_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1971_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1974_inst_ack_0 : boolean;
  signal type_cast_2061_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1974_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1974_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1977_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1977_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1971_inst_req_0 : boolean;
  signal array_obj_ref_2168_index_offset_req_0 : boolean;
  signal RPIPE_Block1_start_1974_inst_req_0 : boolean;
  signal type_cast_2178_inst_ack_0 : boolean;
  signal type_cast_2067_inst_req_0 : boolean;
  signal type_cast_2065_inst_ack_0 : boolean;
  signal type_cast_2273_inst_req_1 : boolean;
  signal type_cast_2178_inst_ack_1 : boolean;
  signal array_obj_ref_2198_index_offset_req_0 : boolean;
  signal type_cast_2273_inst_ack_1 : boolean;
  signal array_obj_ref_2198_index_offset_ack_0 : boolean;
  signal array_obj_ref_2168_index_offset_ack_1 : boolean;
  signal type_cast_2067_inst_ack_0 : boolean;
  signal type_cast_2247_inst_req_0 : boolean;
  signal type_cast_2256_inst_req_1 : boolean;
  signal type_cast_2208_inst_req_0 : boolean;
  signal type_cast_2247_inst_ack_0 : boolean;
  signal ptr_deref_2173_load_0_req_1 : boolean;
  signal type_cast_2208_inst_ack_0 : boolean;
  signal type_cast_2065_inst_req_1 : boolean;
  signal type_cast_2256_inst_ack_1 : boolean;
  signal ptr_deref_2173_load_0_ack_1 : boolean;
  signal type_cast_2065_inst_ack_1 : boolean;
  signal phi_stmt_2062_req_0 : boolean;
  signal array_obj_ref_2198_index_offset_req_1 : boolean;
  signal array_obj_ref_2198_index_offset_ack_1 : boolean;
  signal type_cast_2208_inst_req_1 : boolean;
  signal phi_stmt_2055_req_0 : boolean;
  signal type_cast_2208_inst_ack_1 : boolean;
  signal type_cast_2192_inst_req_0 : boolean;
  signal phi_stmt_2062_req_1 : boolean;
  signal type_cast_2127_inst_req_1 : boolean;
  signal type_cast_2127_inst_ack_0 : boolean;
  signal type_cast_2256_inst_req_0 : boolean;
  signal type_cast_2256_inst_ack_0 : boolean;
  signal addr_of_2169_final_reg_req_0 : boolean;
  signal type_cast_2178_inst_req_0 : boolean;
  signal type_cast_2247_inst_req_1 : boolean;
  signal type_cast_2061_inst_req_1 : boolean;
  signal addr_of_2199_final_reg_req_0 : boolean;
  signal addr_of_2199_final_reg_ack_0 : boolean;
  signal type_cast_2061_inst_ack_1 : boolean;
  signal phi_stmt_2055_req_1 : boolean;
  signal addr_of_2199_final_reg_req_1 : boolean;
  signal phi_stmt_2055_ack_0 : boolean;
  signal type_cast_2127_inst_req_0 : boolean;
  signal if_stmt_2223_branch_req_0 : boolean;
  signal addr_of_2169_final_reg_ack_0 : boolean;
  signal type_cast_2067_inst_req_1 : boolean;
  signal phi_stmt_2062_ack_0 : boolean;
  signal RPIPE_Block1_start_1977_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1977_inst_ack_1 : boolean;
  signal ptr_deref_2202_store_0_ack_1 : boolean;
  signal RPIPE_Block1_start_1980_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1980_inst_ack_0 : boolean;
  signal ptr_deref_2202_store_0_req_1 : boolean;
  signal RPIPE_Block1_start_1980_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1980_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1983_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1983_inst_ack_0 : boolean;
  signal ptr_deref_2173_load_0_ack_0 : boolean;
  signal RPIPE_Block1_start_1983_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1983_inst_ack_1 : boolean;
  signal type_cast_2061_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1986_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1986_inst_ack_0 : boolean;
  signal ptr_deref_2173_load_0_req_0 : boolean;
  signal RPIPE_Block1_start_1986_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1986_inst_ack_1 : boolean;
  signal WPIPE_Block2_done_2288_inst_ack_1 : boolean;
  signal WPIPE_Block2_done_2288_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1989_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1989_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1989_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1989_inst_ack_1 : boolean;
  signal WPIPE_Block2_done_2288_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1992_inst_req_0 : boolean;
  signal ptr_deref_2202_store_0_ack_0 : boolean;
  signal RPIPE_Block1_start_1992_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1992_inst_req_1 : boolean;
  signal ptr_deref_2202_store_0_req_0 : boolean;
  signal RPIPE_Block1_start_1992_inst_ack_1 : boolean;
  signal WPIPE_Block2_done_2288_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1995_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1995_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1995_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1995_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1998_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1998_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1998_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1998_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2001_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2001_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2001_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2001_inst_ack_1 : boolean;
  signal addr_of_2169_final_reg_ack_1 : boolean;
  signal addr_of_2169_final_reg_req_1 : boolean;
  signal if_stmt_2280_branch_ack_0 : boolean;
  signal RPIPE_Block1_start_2004_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2004_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2004_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2004_inst_ack_1 : boolean;
  signal type_cast_2067_inst_ack_1 : boolean;
  signal if_stmt_2280_branch_ack_1 : boolean;
  signal if_stmt_2223_branch_ack_0 : boolean;
  signal type_cast_2015_inst_req_0 : boolean;
  signal type_cast_2015_inst_ack_0 : boolean;
  signal addr_of_2199_final_reg_ack_1 : boolean;
  signal type_cast_2273_inst_ack_0 : boolean;
  signal type_cast_2015_inst_req_1 : boolean;
  signal type_cast_2015_inst_ack_1 : boolean;
  signal type_cast_2192_inst_ack_1 : boolean;
  signal type_cast_2273_inst_req_0 : boolean;
  signal type_cast_2019_inst_req_0 : boolean;
  signal type_cast_2019_inst_ack_0 : boolean;
  signal type_cast_2019_inst_req_1 : boolean;
  signal type_cast_2019_inst_ack_1 : boolean;
  signal if_stmt_2223_branch_ack_1 : boolean;
  signal type_cast_2192_inst_req_1 : boolean;
  signal type_cast_2029_inst_req_0 : boolean;
  signal type_cast_2029_inst_ack_0 : boolean;
  signal type_cast_2029_inst_req_1 : boolean;
  signal type_cast_2029_inst_ack_1 : boolean;
  signal if_stmt_2280_branch_req_0 : boolean;
  signal type_cast_2247_inst_ack_1 : boolean;
  signal type_cast_2192_inst_ack_0 : boolean;
  signal type_cast_2148_inst_req_0 : boolean;
  signal type_cast_2148_inst_ack_0 : boolean;
  signal type_cast_2148_inst_req_1 : boolean;
  signal type_cast_2148_inst_ack_1 : boolean;
  signal type_cast_2162_inst_req_0 : boolean;
  signal type_cast_2162_inst_ack_0 : boolean;
  signal type_cast_2162_inst_req_1 : boolean;
  signal type_cast_2162_inst_ack_1 : boolean;
  signal type_cast_2127_inst_ack_1 : boolean;
  signal phi_stmt_2121_req_1 : boolean;
  signal phi_stmt_2121_req_0 : boolean;
  signal phi_stmt_2121_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeC_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeC_CP_4929_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeC_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_4929_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeC_CP_4929_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_4929_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeC_CP_4929: Block -- control-path 
    signal convTransposeC_CP_4929_elements: BooleanArray(89 downto 0);
    -- 
  begin -- 
    convTransposeC_CP_4929_elements(0) <= convTransposeC_CP_4929_start;
    convTransposeC_CP_4929_symbol <= convTransposeC_CP_4929_elements(67);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1971_sample_start_
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1969/branch_block_stmt_1969__entry__
      -- CP-element group 0: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/$entry
      -- CP-element group 0: 	 branch_block_stmt_1969/$entry
      -- CP-element group 0: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005__entry__
      -- CP-element group 0: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1971_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1971_Sample/rr
      -- 
    rr_4977_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4977_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(0), ack => RPIPE_Block1_start_1971_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1971_update_start_
      -- CP-element group 1: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1971_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1971_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1971_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1971_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1971_Update/$entry
      -- 
    ra_4978_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1971_inst_ack_0, ack => convTransposeC_CP_4929_elements(1)); -- 
    cr_4982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(1), ack => RPIPE_Block1_start_1971_inst_req_1); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1971_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1971_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1974_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1971_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1974_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1974_Sample/rr
      -- 
    ca_4983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1971_inst_ack_1, ack => convTransposeC_CP_4929_elements(2)); -- 
    rr_4991_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4991_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(2), ack => RPIPE_Block1_start_1974_inst_req_0); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1974_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1974_Update/cr
      -- CP-element group 3: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1974_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1974_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1974_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1974_update_start_
      -- 
    ra_4992_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1974_inst_ack_0, ack => convTransposeC_CP_4929_elements(3)); -- 
    cr_4996_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4996_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(3), ack => RPIPE_Block1_start_1974_inst_req_1); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1974_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1977_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1974_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1977_Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1974_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1977_Sample/$entry
      -- 
    ca_4997_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1974_inst_ack_1, ack => convTransposeC_CP_4929_elements(4)); -- 
    rr_5005_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5005_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(4), ack => RPIPE_Block1_start_1977_inst_req_0); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1977_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1977_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1977_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1977_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1977_update_start_
      -- CP-element group 5: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1977_Update/cr
      -- 
    ra_5006_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1977_inst_ack_0, ack => convTransposeC_CP_4929_elements(5)); -- 
    cr_5010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(5), ack => RPIPE_Block1_start_1977_inst_req_1); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1977_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1977_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1977_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1980_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1980_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1980_Sample/rr
      -- 
    ca_5011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1977_inst_ack_1, ack => convTransposeC_CP_4929_elements(6)); -- 
    rr_5019_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5019_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(6), ack => RPIPE_Block1_start_1980_inst_req_0); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1980_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1980_update_start_
      -- CP-element group 7: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1980_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1980_Sample/ra
      -- CP-element group 7: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1980_Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1980_Update/cr
      -- 
    ra_5020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1980_inst_ack_0, ack => convTransposeC_CP_4929_elements(7)); -- 
    cr_5024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(7), ack => RPIPE_Block1_start_1980_inst_req_1); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1980_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1980_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1980_Update/ca
      -- CP-element group 8: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1983_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1983_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1983_Sample/rr
      -- 
    ca_5025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1980_inst_ack_1, ack => convTransposeC_CP_4929_elements(8)); -- 
    rr_5033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(8), ack => RPIPE_Block1_start_1983_inst_req_0); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1983_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1983_update_start_
      -- CP-element group 9: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1983_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1983_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1983_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1983_Update/cr
      -- 
    ra_5034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1983_inst_ack_0, ack => convTransposeC_CP_4929_elements(9)); -- 
    cr_5038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(9), ack => RPIPE_Block1_start_1983_inst_req_1); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1983_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1983_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1983_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1986_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1986_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1986_Sample/rr
      -- 
    ca_5039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1983_inst_ack_1, ack => convTransposeC_CP_4929_elements(10)); -- 
    rr_5047_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5047_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(10), ack => RPIPE_Block1_start_1986_inst_req_0); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1986_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1986_update_start_
      -- CP-element group 11: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1986_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1986_Sample/ra
      -- CP-element group 11: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1986_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1986_Update/cr
      -- 
    ra_5048_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1986_inst_ack_0, ack => convTransposeC_CP_4929_elements(11)); -- 
    cr_5052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(11), ack => RPIPE_Block1_start_1986_inst_req_1); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1986_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1986_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1986_Update/ca
      -- CP-element group 12: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1989_sample_start_
      -- CP-element group 12: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1989_Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1989_Sample/rr
      -- 
    ca_5053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1986_inst_ack_1, ack => convTransposeC_CP_4929_elements(12)); -- 
    rr_5061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(12), ack => RPIPE_Block1_start_1989_inst_req_0); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1989_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1989_update_start_
      -- CP-element group 13: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1989_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1989_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1989_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1989_Update/cr
      -- 
    ra_5062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1989_inst_ack_0, ack => convTransposeC_CP_4929_elements(13)); -- 
    cr_5066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(13), ack => RPIPE_Block1_start_1989_inst_req_1); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1989_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1989_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1989_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1992_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1992_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1992_Sample/rr
      -- 
    ca_5067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1989_inst_ack_1, ack => convTransposeC_CP_4929_elements(14)); -- 
    rr_5075_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5075_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(14), ack => RPIPE_Block1_start_1992_inst_req_0); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1992_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1992_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1992_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1992_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1992_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1992_Update/cr
      -- 
    ra_5076_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1992_inst_ack_0, ack => convTransposeC_CP_4929_elements(15)); -- 
    cr_5080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(15), ack => RPIPE_Block1_start_1992_inst_req_1); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1992_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1992_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1992_Update/ca
      -- CP-element group 16: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1995_sample_start_
      -- CP-element group 16: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1995_Sample/$entry
      -- CP-element group 16: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1995_Sample/rr
      -- 
    ca_5081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1992_inst_ack_1, ack => convTransposeC_CP_4929_elements(16)); -- 
    rr_5089_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5089_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(16), ack => RPIPE_Block1_start_1995_inst_req_0); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1995_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1995_update_start_
      -- CP-element group 17: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1995_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1995_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1995_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1995_Update/cr
      -- 
    ra_5090_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1995_inst_ack_0, ack => convTransposeC_CP_4929_elements(17)); -- 
    cr_5094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(17), ack => RPIPE_Block1_start_1995_inst_req_1); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1995_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1995_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1995_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1998_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1998_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1998_Sample/rr
      -- 
    ca_5095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1995_inst_ack_1, ack => convTransposeC_CP_4929_elements(18)); -- 
    rr_5103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(18), ack => RPIPE_Block1_start_1998_inst_req_0); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1998_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1998_update_start_
      -- CP-element group 19: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1998_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1998_Sample/ra
      -- CP-element group 19: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1998_Update/$entry
      -- CP-element group 19: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1998_Update/cr
      -- 
    ra_5104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1998_inst_ack_0, ack => convTransposeC_CP_4929_elements(19)); -- 
    cr_5108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(19), ack => RPIPE_Block1_start_1998_inst_req_1); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1998_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1998_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_1998_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_2001_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_2001_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_2001_Sample/rr
      -- 
    ca_5109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1998_inst_ack_1, ack => convTransposeC_CP_4929_elements(20)); -- 
    rr_5117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(20), ack => RPIPE_Block1_start_2001_inst_req_0); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_2001_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_2001_update_start_
      -- CP-element group 21: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_2001_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_2001_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_2001_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_2001_Update/cr
      -- 
    ra_5118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2001_inst_ack_0, ack => convTransposeC_CP_4929_elements(21)); -- 
    cr_5122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(21), ack => RPIPE_Block1_start_2001_inst_req_1); -- 
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (6) 
      -- CP-element group 22: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_2001_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_2001_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_2001_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_2004_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_2004_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_2004_Sample/rr
      -- 
    ca_5123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2001_inst_ack_1, ack => convTransposeC_CP_4929_elements(22)); -- 
    rr_5131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(22), ack => RPIPE_Block1_start_2004_inst_req_0); -- 
    -- CP-element group 23:  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (6) 
      -- CP-element group 23: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_2004_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_2004_update_start_
      -- CP-element group 23: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_2004_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_2004_Sample/ra
      -- CP-element group 23: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_2004_Update/$entry
      -- CP-element group 23: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_2004_Update/cr
      -- 
    ra_5132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2004_inst_ack_0, ack => convTransposeC_CP_4929_elements(23)); -- 
    cr_5136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(23), ack => RPIPE_Block1_start_2004_inst_req_1); -- 
    -- CP-element group 24:  fork  transition  place  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24: 	26 
    -- CP-element group 24: 	27 
    -- CP-element group 24: 	28 
    -- CP-element group 24: 	29 
    -- CP-element group 24: 	30 
    -- CP-element group 24:  members (25) 
      -- CP-element group 24: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/$exit
      -- CP-element group 24: 	 branch_block_stmt_1969/assign_stmt_2012_to_assign_stmt_2052__entry__
      -- CP-element group 24: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005__exit__
      -- CP-element group 24: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_2004_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_2004_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_1969/assign_stmt_1972_to_assign_stmt_2005/RPIPE_Block1_start_2004_Update/ca
      -- CP-element group 24: 	 branch_block_stmt_1969/assign_stmt_2012_to_assign_stmt_2052/$entry
      -- CP-element group 24: 	 branch_block_stmt_1969/assign_stmt_2012_to_assign_stmt_2052/type_cast_2015_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1969/assign_stmt_2012_to_assign_stmt_2052/type_cast_2015_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1969/assign_stmt_2012_to_assign_stmt_2052/type_cast_2015_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_1969/assign_stmt_2012_to_assign_stmt_2052/type_cast_2015_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_1969/assign_stmt_2012_to_assign_stmt_2052/type_cast_2015_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1969/assign_stmt_2012_to_assign_stmt_2052/type_cast_2015_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_1969/assign_stmt_2012_to_assign_stmt_2052/type_cast_2019_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1969/assign_stmt_2012_to_assign_stmt_2052/type_cast_2019_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1969/assign_stmt_2012_to_assign_stmt_2052/type_cast_2019_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_1969/assign_stmt_2012_to_assign_stmt_2052/type_cast_2019_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_1969/assign_stmt_2012_to_assign_stmt_2052/type_cast_2019_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1969/assign_stmt_2012_to_assign_stmt_2052/type_cast_2019_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_1969/assign_stmt_2012_to_assign_stmt_2052/type_cast_2029_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1969/assign_stmt_2012_to_assign_stmt_2052/type_cast_2029_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1969/assign_stmt_2012_to_assign_stmt_2052/type_cast_2029_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_1969/assign_stmt_2012_to_assign_stmt_2052/type_cast_2029_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_1969/assign_stmt_2012_to_assign_stmt_2052/type_cast_2029_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1969/assign_stmt_2012_to_assign_stmt_2052/type_cast_2029_Update/cr
      -- 
    ca_5137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2004_inst_ack_1, ack => convTransposeC_CP_4929_elements(24)); -- 
    rr_5148_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5148_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(24), ack => type_cast_2015_inst_req_0); -- 
    cr_5153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(24), ack => type_cast_2015_inst_req_1); -- 
    rr_5162_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5162_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(24), ack => type_cast_2019_inst_req_0); -- 
    cr_5167_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5167_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(24), ack => type_cast_2019_inst_req_1); -- 
    rr_5176_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5176_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(24), ack => type_cast_2029_inst_req_0); -- 
    cr_5181_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5181_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(24), ack => type_cast_2029_inst_req_1); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_1969/assign_stmt_2012_to_assign_stmt_2052/type_cast_2015_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_1969/assign_stmt_2012_to_assign_stmt_2052/type_cast_2015_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_1969/assign_stmt_2012_to_assign_stmt_2052/type_cast_2015_Sample/ra
      -- 
    ra_5149_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2015_inst_ack_0, ack => convTransposeC_CP_4929_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	31 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1969/assign_stmt_2012_to_assign_stmt_2052/type_cast_2015_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_1969/assign_stmt_2012_to_assign_stmt_2052/type_cast_2015_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_1969/assign_stmt_2012_to_assign_stmt_2052/type_cast_2015_Update/ca
      -- 
    ca_5154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2015_inst_ack_1, ack => convTransposeC_CP_4929_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	24 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1969/assign_stmt_2012_to_assign_stmt_2052/type_cast_2019_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_1969/assign_stmt_2012_to_assign_stmt_2052/type_cast_2019_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_1969/assign_stmt_2012_to_assign_stmt_2052/type_cast_2019_Sample/ra
      -- 
    ra_5163_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2019_inst_ack_0, ack => convTransposeC_CP_4929_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	24 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	31 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1969/assign_stmt_2012_to_assign_stmt_2052/type_cast_2019_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_1969/assign_stmt_2012_to_assign_stmt_2052/type_cast_2019_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_1969/assign_stmt_2012_to_assign_stmt_2052/type_cast_2019_Update/ca
      -- 
    ca_5168_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2019_inst_ack_1, ack => convTransposeC_CP_4929_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	24 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_1969/assign_stmt_2012_to_assign_stmt_2052/type_cast_2029_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_1969/assign_stmt_2012_to_assign_stmt_2052/type_cast_2029_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_1969/assign_stmt_2012_to_assign_stmt_2052/type_cast_2029_Sample/ra
      -- 
    ra_5177_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2029_inst_ack_0, ack => convTransposeC_CP_4929_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	24 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1969/assign_stmt_2012_to_assign_stmt_2052/type_cast_2029_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_1969/assign_stmt_2012_to_assign_stmt_2052/type_cast_2029_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_1969/assign_stmt_2012_to_assign_stmt_2052/type_cast_2029_Update/ca
      -- 
    ca_5182_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2029_inst_ack_1, ack => convTransposeC_CP_4929_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  place  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	26 
    -- CP-element group 31: 	28 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	68 
    -- CP-element group 31: 	69 
    -- CP-element group 31: 	71 
    -- CP-element group 31:  members (14) 
      -- CP-element group 31: 	 branch_block_stmt_1969/assign_stmt_2012_to_assign_stmt_2052__exit__
      -- CP-element group 31: 	 branch_block_stmt_1969/entry_whilex_xbodyx_xouter
      -- CP-element group 31: 	 branch_block_stmt_1969/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/type_cast_2065/SplitProtocol/Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_1969/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/type_cast_2065/SplitProtocol/$entry
      -- CP-element group 31: 	 branch_block_stmt_1969/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/type_cast_2065/SplitProtocol/Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1969/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/type_cast_2065/$entry
      -- CP-element group 31: 	 branch_block_stmt_1969/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/type_cast_2065/SplitProtocol/Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_1969/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/type_cast_2065/SplitProtocol/Update/cr
      -- CP-element group 31: 	 branch_block_stmt_1969/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2055/$entry
      -- CP-element group 31: 	 branch_block_stmt_1969/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/$entry
      -- CP-element group 31: 	 branch_block_stmt_1969/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/$entry
      -- CP-element group 31: 	 branch_block_stmt_1969/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2062/$entry
      -- CP-element group 31: 	 branch_block_stmt_1969/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 31: 	 branch_block_stmt_1969/assign_stmt_2012_to_assign_stmt_2052/$exit
      -- 
    rr_5572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(31), ack => type_cast_2065_inst_req_0); -- 
    cr_5577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(31), ack => type_cast_2065_inst_req_1); -- 
    convTransposeC_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_4929_elements(26) & convTransposeC_CP_4929_elements(28) & convTransposeC_CP_4929_elements(30);
      gj_convTransposeC_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_4929_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	89 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2148_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2148_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2148_Sample/ra
      -- 
    ra_5197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2148_inst_ack_0, ack => convTransposeC_CP_4929_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	89 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2148_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2148_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2148_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2162_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2162_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2162_Sample/rr
      -- 
    ca_5202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2148_inst_ack_1, ack => convTransposeC_CP_4929_elements(33)); -- 
    rr_5210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(33), ack => type_cast_2162_inst_req_0); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2162_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2162_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2162_Sample/ra
      -- 
    ra_5211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2162_inst_ack_0, ack => convTransposeC_CP_4929_elements(34)); -- 
    -- CP-element group 35:  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	89 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (16) 
      -- CP-element group 35: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2168_final_index_sum_regn_Sample/req
      -- CP-element group 35: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2168_final_index_sum_regn_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2162_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2162_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2162_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2168_index_resized_1
      -- CP-element group 35: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2168_index_scaled_1
      -- CP-element group 35: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2168_index_computed_1
      -- CP-element group 35: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2168_index_resize_1/$entry
      -- CP-element group 35: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2168_index_resize_1/$exit
      -- CP-element group 35: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2168_index_resize_1/index_resize_req
      -- CP-element group 35: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2168_index_resize_1/index_resize_ack
      -- CP-element group 35: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2168_index_scale_1/$entry
      -- CP-element group 35: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2168_index_scale_1/$exit
      -- CP-element group 35: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2168_index_scale_1/scale_rename_req
      -- CP-element group 35: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2168_index_scale_1/scale_rename_ack
      -- 
    ca_5216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2162_inst_ack_1, ack => convTransposeC_CP_4929_elements(35)); -- 
    req_5241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(35), ack => array_obj_ref_2168_index_offset_req_0); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	55 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2168_final_index_sum_regn_Sample/ack
      -- CP-element group 36: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2168_final_index_sum_regn_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2168_final_index_sum_regn_sample_complete
      -- 
    ack_5242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2168_index_offset_ack_0, ack => convTransposeC_CP_4929_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	89 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (11) 
      -- CP-element group 37: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2168_final_index_sum_regn_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2168_final_index_sum_regn_Update/ack
      -- CP-element group 37: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2168_base_plus_offset/$entry
      -- CP-element group 37: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2168_base_plus_offset/$exit
      -- CP-element group 37: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2168_base_plus_offset/sum_rename_req
      -- CP-element group 37: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2168_base_plus_offset/sum_rename_ack
      -- CP-element group 37: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/addr_of_2169_request/$entry
      -- CP-element group 37: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/addr_of_2169_request/req
      -- CP-element group 37: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/addr_of_2169_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2168_root_address_calculated
      -- CP-element group 37: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2168_offset_calculated
      -- 
    ack_5247_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2168_index_offset_ack_1, ack => convTransposeC_CP_4929_elements(37)); -- 
    req_5256_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5256_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(37), ack => addr_of_2169_final_reg_req_0); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/addr_of_2169_request/$exit
      -- CP-element group 38: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/addr_of_2169_request/ack
      -- CP-element group 38: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/addr_of_2169_sample_completed_
      -- 
    ack_5257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2169_final_reg_ack_0, ack => convTransposeC_CP_4929_elements(38)); -- 
    -- CP-element group 39:  join  fork  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	89 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (24) 
      -- CP-element group 39: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2173_base_addr_resize/base_resize_ack
      -- CP-element group 39: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2173_base_addr_resize/base_resize_req
      -- CP-element group 39: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2173_word_addrgen/$entry
      -- CP-element group 39: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/addr_of_2169_complete/$exit
      -- CP-element group 39: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2173_base_plus_offset/$entry
      -- CP-element group 39: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2173_base_plus_offset/$exit
      -- CP-element group 39: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2173_base_plus_offset/sum_rename_req
      -- CP-element group 39: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2173_base_plus_offset/sum_rename_ack
      -- CP-element group 39: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2173_base_addr_resize/$exit
      -- CP-element group 39: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2173_base_addr_resize/$entry
      -- CP-element group 39: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2173_base_address_resized
      -- CP-element group 39: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2173_root_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2173_word_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2173_base_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2173_Sample/word_access_start/word_0/rr
      -- CP-element group 39: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2173_Sample/word_access_start/word_0/$entry
      -- CP-element group 39: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2173_Sample/word_access_start/$entry
      -- CP-element group 39: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2173_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/addr_of_2169_complete/ack
      -- CP-element group 39: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2173_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2173_word_addrgen/root_register_ack
      -- CP-element group 39: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2173_word_addrgen/root_register_req
      -- CP-element group 39: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2173_word_addrgen/$exit
      -- CP-element group 39: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/addr_of_2169_update_completed_
      -- 
    ack_5262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2169_final_reg_ack_1, ack => convTransposeC_CP_4929_elements(39)); -- 
    rr_5295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(39), ack => ptr_deref_2173_load_0_req_0); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (5) 
      -- CP-element group 40: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2173_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2173_Sample/word_access_start/word_0/ra
      -- CP-element group 40: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2173_Sample/word_access_start/word_0/$exit
      -- CP-element group 40: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2173_Sample/word_access_start/$exit
      -- CP-element group 40: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2173_Sample/$exit
      -- 
    ra_5296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2173_load_0_ack_0, ack => convTransposeC_CP_4929_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	89 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	50 
    -- CP-element group 41:  members (9) 
      -- CP-element group 41: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2173_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2173_Update/word_access_complete/$exit
      -- CP-element group 41: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2173_Update/word_access_complete/word_0/$exit
      -- CP-element group 41: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2173_Update/word_access_complete/word_0/ca
      -- CP-element group 41: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2173_Update/ptr_deref_2173_Merge/$entry
      -- CP-element group 41: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2173_Update/ptr_deref_2173_Merge/$exit
      -- CP-element group 41: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2173_Update/ptr_deref_2173_Merge/merge_req
      -- CP-element group 41: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2173_Update/ptr_deref_2173_Merge/merge_ack
      -- CP-element group 41: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2173_update_completed_
      -- 
    ca_5307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2173_load_0_ack_1, ack => convTransposeC_CP_4929_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	89 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2178_Sample/ra
      -- CP-element group 42: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2178_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2178_Sample/$exit
      -- 
    ra_5321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2178_inst_ack_0, ack => convTransposeC_CP_4929_elements(42)); -- 
    -- CP-element group 43:  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	89 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (6) 
      -- CP-element group 43: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2178_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2178_Update/ca
      -- CP-element group 43: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2192_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2178_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2192_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2192_Sample/rr
      -- 
    ca_5326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2178_inst_ack_1, ack => convTransposeC_CP_4929_elements(43)); -- 
    rr_5334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(43), ack => type_cast_2192_inst_req_0); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2192_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2192_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2192_Sample/ra
      -- 
    ra_5335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2192_inst_ack_0, ack => convTransposeC_CP_4929_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	89 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (16) 
      -- CP-element group 45: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2198_index_scale_1/scale_rename_ack
      -- CP-element group 45: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2198_index_scale_1/scale_rename_req
      -- CP-element group 45: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2198_final_index_sum_regn_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2198_final_index_sum_regn_Sample/req
      -- CP-element group 45: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2192_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2198_index_scale_1/$exit
      -- CP-element group 45: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2198_index_scale_1/$entry
      -- CP-element group 45: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2198_index_resize_1/index_resize_ack
      -- CP-element group 45: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2198_index_resize_1/index_resize_req
      -- CP-element group 45: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2198_index_resize_1/$exit
      -- CP-element group 45: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2198_index_resize_1/$entry
      -- CP-element group 45: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2198_index_computed_1
      -- CP-element group 45: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2198_index_scaled_1
      -- CP-element group 45: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2198_index_resized_1
      -- CP-element group 45: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2192_Update/ca
      -- CP-element group 45: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2192_Update/$exit
      -- 
    ca_5340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2192_inst_ack_1, ack => convTransposeC_CP_4929_elements(45)); -- 
    req_5365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(45), ack => array_obj_ref_2198_index_offset_req_0); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	55 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2198_final_index_sum_regn_sample_complete
      -- CP-element group 46: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2198_final_index_sum_regn_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2198_final_index_sum_regn_Sample/ack
      -- 
    ack_5366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2198_index_offset_ack_0, ack => convTransposeC_CP_4929_elements(46)); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	89 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (11) 
      -- CP-element group 47: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2198_final_index_sum_regn_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2198_final_index_sum_regn_Update/ack
      -- CP-element group 47: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2198_base_plus_offset/$entry
      -- CP-element group 47: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2198_base_plus_offset/$exit
      -- CP-element group 47: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2198_base_plus_offset/sum_rename_req
      -- CP-element group 47: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2198_base_plus_offset/sum_rename_ack
      -- CP-element group 47: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/addr_of_2199_request/$entry
      -- CP-element group 47: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/addr_of_2199_request/req
      -- CP-element group 47: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2198_offset_calculated
      -- CP-element group 47: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2198_root_address_calculated
      -- CP-element group 47: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/addr_of_2199_sample_start_
      -- 
    ack_5371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2198_index_offset_ack_1, ack => convTransposeC_CP_4929_elements(47)); -- 
    req_5380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(47), ack => addr_of_2199_final_reg_req_0); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/addr_of_2199_request/$exit
      -- CP-element group 48: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/addr_of_2199_request/ack
      -- CP-element group 48: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/addr_of_2199_sample_completed_
      -- 
    ack_5381_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2199_final_reg_ack_0, ack => convTransposeC_CP_4929_elements(48)); -- 
    -- CP-element group 49:  fork  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	89 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (19) 
      -- CP-element group 49: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2202_base_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2202_word_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2202_root_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2202_base_address_resized
      -- CP-element group 49: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2202_base_addr_resize/$entry
      -- CP-element group 49: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2202_base_addr_resize/$exit
      -- CP-element group 49: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2202_base_addr_resize/base_resize_req
      -- CP-element group 49: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2202_base_addr_resize/base_resize_ack
      -- CP-element group 49: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2202_base_plus_offset/$entry
      -- CP-element group 49: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2202_base_plus_offset/$exit
      -- CP-element group 49: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2202_base_plus_offset/sum_rename_req
      -- CP-element group 49: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2202_base_plus_offset/sum_rename_ack
      -- CP-element group 49: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/addr_of_2199_complete/$exit
      -- CP-element group 49: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/addr_of_2199_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/addr_of_2199_complete/ack
      -- CP-element group 49: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2202_word_addrgen/root_register_ack
      -- CP-element group 49: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2202_word_addrgen/root_register_req
      -- CP-element group 49: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2202_word_addrgen/$exit
      -- CP-element group 49: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2202_word_addrgen/$entry
      -- 
    ack_5386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2199_final_reg_ack_1, ack => convTransposeC_CP_4929_elements(49)); -- 
    -- CP-element group 50:  join  transition  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	41 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2202_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2202_Sample/word_access_start/word_0/rr
      -- CP-element group 50: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2202_Sample/word_access_start/word_0/$entry
      -- CP-element group 50: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2202_Sample/word_access_start/$entry
      -- CP-element group 50: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2202_Sample/ptr_deref_2202_Split/split_ack
      -- CP-element group 50: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2202_Sample/ptr_deref_2202_Split/split_req
      -- CP-element group 50: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2202_Sample/ptr_deref_2202_Split/$exit
      -- CP-element group 50: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2202_Sample/ptr_deref_2202_Split/$entry
      -- CP-element group 50: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2202_Sample/$entry
      -- 
    rr_5424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(50), ack => ptr_deref_2202_store_0_req_0); -- 
    convTransposeC_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_4929_elements(41) & convTransposeC_CP_4929_elements(49);
      gj_convTransposeC_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_4929_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (5) 
      -- CP-element group 51: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2202_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2202_Sample/word_access_start/word_0/ra
      -- CP-element group 51: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2202_Sample/word_access_start/word_0/$exit
      -- CP-element group 51: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2202_Sample/word_access_start/$exit
      -- CP-element group 51: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2202_Sample/$exit
      -- 
    ra_5425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2202_store_0_ack_0, ack => convTransposeC_CP_4929_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	89 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	55 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2202_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2202_Update/word_access_complete/word_0/ca
      -- CP-element group 52: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2202_Update/word_access_complete/word_0/$exit
      -- CP-element group 52: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2202_Update/word_access_complete/$exit
      -- CP-element group 52: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2202_Update/$exit
      -- 
    ca_5436_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2202_store_0_ack_1, ack => convTransposeC_CP_4929_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	89 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2208_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2208_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2208_Sample/ra
      -- 
    ra_5445_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2208_inst_ack_0, ack => convTransposeC_CP_4929_elements(53)); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	89 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2208_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2208_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2208_Update/ca
      -- 
    ca_5450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2208_inst_ack_1, ack => convTransposeC_CP_4929_elements(54)); -- 
    -- CP-element group 55:  branch  join  transition  place  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	36 
    -- CP-element group 55: 	46 
    -- CP-element group 55: 	52 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (10) 
      -- CP-element group 55: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222__exit__
      -- CP-element group 55: 	 branch_block_stmt_1969/if_stmt_2223__entry__
      -- CP-element group 55: 	 branch_block_stmt_1969/if_stmt_2223_dead_link/$entry
      -- CP-element group 55: 	 branch_block_stmt_1969/if_stmt_2223_eval_test/$entry
      -- CP-element group 55: 	 branch_block_stmt_1969/if_stmt_2223_eval_test/$exit
      -- CP-element group 55: 	 branch_block_stmt_1969/if_stmt_2223_eval_test/branch_req
      -- CP-element group 55: 	 branch_block_stmt_1969/if_stmt_2223_else_link/$entry
      -- CP-element group 55: 	 branch_block_stmt_1969/if_stmt_2223_if_link/$entry
      -- CP-element group 55: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/$exit
      -- CP-element group 55: 	 branch_block_stmt_1969/R_cmp_2224_place
      -- 
    branch_req_5458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(55), ack => if_stmt_2223_branch_req_0); -- 
    convTransposeC_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_4929_elements(36) & convTransposeC_CP_4929_elements(46) & convTransposeC_CP_4929_elements(52) & convTransposeC_CP_4929_elements(54);
      gj_convTransposeC_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_4929_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	84 
    -- CP-element group 56: 	85 
    -- CP-element group 56:  members (24) 
      -- CP-element group 56: 	 branch_block_stmt_1969/ifx_xthen_whilex_xbody
      -- CP-element group 56: 	 branch_block_stmt_1969/merge_stmt_2229_PhiReqMerge
      -- CP-element group 56: 	 branch_block_stmt_1969/merge_stmt_2229__exit__
      -- CP-element group 56: 	 branch_block_stmt_1969/assign_stmt_2235__entry__
      -- CP-element group 56: 	 branch_block_stmt_1969/assign_stmt_2235__exit__
      -- CP-element group 56: 	 branch_block_stmt_1969/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2121/phi_stmt_2121_sources/type_cast_2127/SplitProtocol/Update/cr
      -- CP-element group 56: 	 branch_block_stmt_1969/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2121/$entry
      -- CP-element group 56: 	 branch_block_stmt_1969/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2121/phi_stmt_2121_sources/$entry
      -- CP-element group 56: 	 branch_block_stmt_1969/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2121/phi_stmt_2121_sources/type_cast_2127/SplitProtocol/$entry
      -- CP-element group 56: 	 branch_block_stmt_1969/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2121/phi_stmt_2121_sources/type_cast_2127/SplitProtocol/Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_1969/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2121/phi_stmt_2121_sources/type_cast_2127/$entry
      -- CP-element group 56: 	 branch_block_stmt_1969/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 56: 	 branch_block_stmt_1969/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2121/phi_stmt_2121_sources/type_cast_2127/SplitProtocol/Sample/rr
      -- CP-element group 56: 	 branch_block_stmt_1969/assign_stmt_2235/$exit
      -- CP-element group 56: 	 branch_block_stmt_1969/assign_stmt_2235/$entry
      -- CP-element group 56: 	 branch_block_stmt_1969/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2121/phi_stmt_2121_sources/type_cast_2127/SplitProtocol/Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_1969/if_stmt_2223_if_link/if_choice_transition
      -- CP-element group 56: 	 branch_block_stmt_1969/if_stmt_2223_if_link/$exit
      -- CP-element group 56: 	 branch_block_stmt_1969/whilex_xbody_ifx_xthen
      -- CP-element group 56: 	 branch_block_stmt_1969/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 56: 	 branch_block_stmt_1969/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 56: 	 branch_block_stmt_1969/merge_stmt_2229_PhiAck/$entry
      -- CP-element group 56: 	 branch_block_stmt_1969/merge_stmt_2229_PhiAck/$exit
      -- CP-element group 56: 	 branch_block_stmt_1969/merge_stmt_2229_PhiAck/dummy
      -- 
    if_choice_transition_5463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2223_branch_ack_1, ack => convTransposeC_CP_4929_elements(56)); -- 
    cr_5666_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5666_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(56), ack => type_cast_2127_inst_req_1); -- 
    rr_5661_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5661_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(56), ack => type_cast_2127_inst_req_0); -- 
    -- CP-element group 57:  fork  transition  place  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57: 	59 
    -- CP-element group 57: 	61 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (24) 
      -- CP-element group 57: 	 branch_block_stmt_1969/merge_stmt_2237__exit__
      -- CP-element group 57: 	 branch_block_stmt_1969/assign_stmt_2243_to_assign_stmt_2279__entry__
      -- CP-element group 57: 	 branch_block_stmt_1969/assign_stmt_2243_to_assign_stmt_2279/type_cast_2247_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_1969/assign_stmt_2243_to_assign_stmt_2279/type_cast_2273_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_1969/merge_stmt_2237_PhiReqMerge
      -- CP-element group 57: 	 branch_block_stmt_1969/assign_stmt_2243_to_assign_stmt_2279/type_cast_2247_Sample/rr
      -- CP-element group 57: 	 branch_block_stmt_1969/assign_stmt_2243_to_assign_stmt_2279/type_cast_2256_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_1969/assign_stmt_2243_to_assign_stmt_2279/type_cast_2247_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_1969/assign_stmt_2243_to_assign_stmt_2279/type_cast_2247_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_1969/assign_stmt_2243_to_assign_stmt_2279/type_cast_2273_update_start_
      -- CP-element group 57: 	 branch_block_stmt_1969/assign_stmt_2243_to_assign_stmt_2279/type_cast_2247_update_start_
      -- CP-element group 57: 	 branch_block_stmt_1969/assign_stmt_2243_to_assign_stmt_2279/type_cast_2247_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_1969/assign_stmt_2243_to_assign_stmt_2279/$entry
      -- CP-element group 57: 	 branch_block_stmt_1969/assign_stmt_2243_to_assign_stmt_2279/type_cast_2256_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_1969/if_stmt_2223_else_link/else_choice_transition
      -- CP-element group 57: 	 branch_block_stmt_1969/assign_stmt_2243_to_assign_stmt_2279/type_cast_2273_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_1969/if_stmt_2223_else_link/$exit
      -- CP-element group 57: 	 branch_block_stmt_1969/assign_stmt_2243_to_assign_stmt_2279/type_cast_2256_update_start_
      -- CP-element group 57: 	 branch_block_stmt_1969/whilex_xbody_ifx_xelse
      -- CP-element group 57: 	 branch_block_stmt_1969/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 57: 	 branch_block_stmt_1969/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 57: 	 branch_block_stmt_1969/merge_stmt_2237_PhiAck/$entry
      -- CP-element group 57: 	 branch_block_stmt_1969/merge_stmt_2237_PhiAck/$exit
      -- CP-element group 57: 	 branch_block_stmt_1969/merge_stmt_2237_PhiAck/dummy
      -- 
    else_choice_transition_5467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2223_branch_ack_0, ack => convTransposeC_CP_4929_elements(57)); -- 
    cr_5516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(57), ack => type_cast_2273_inst_req_1); -- 
    rr_5483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(57), ack => type_cast_2247_inst_req_0); -- 
    cr_5502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(57), ack => type_cast_2256_inst_req_1); -- 
    cr_5488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(57), ack => type_cast_2247_inst_req_1); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_1969/assign_stmt_2243_to_assign_stmt_2279/type_cast_2247_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_1969/assign_stmt_2243_to_assign_stmt_2279/type_cast_2247_Sample/ra
      -- CP-element group 58: 	 branch_block_stmt_1969/assign_stmt_2243_to_assign_stmt_2279/type_cast_2247_sample_completed_
      -- 
    ra_5484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2247_inst_ack_0, ack => convTransposeC_CP_4929_elements(58)); -- 
    -- CP-element group 59:  transition  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (6) 
      -- CP-element group 59: 	 branch_block_stmt_1969/assign_stmt_2243_to_assign_stmt_2279/type_cast_2247_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_1969/assign_stmt_2243_to_assign_stmt_2279/type_cast_2256_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_1969/assign_stmt_2243_to_assign_stmt_2279/type_cast_2247_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_1969/assign_stmt_2243_to_assign_stmt_2279/type_cast_2256_Sample/rr
      -- CP-element group 59: 	 branch_block_stmt_1969/assign_stmt_2243_to_assign_stmt_2279/type_cast_2256_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_1969/assign_stmt_2243_to_assign_stmt_2279/type_cast_2247_Update/ca
      -- 
    ca_5489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2247_inst_ack_1, ack => convTransposeC_CP_4929_elements(59)); -- 
    rr_5497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(59), ack => type_cast_2256_inst_req_0); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_1969/assign_stmt_2243_to_assign_stmt_2279/type_cast_2256_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_1969/assign_stmt_2243_to_assign_stmt_2279/type_cast_2256_Sample/ra
      -- CP-element group 60: 	 branch_block_stmt_1969/assign_stmt_2243_to_assign_stmt_2279/type_cast_2256_sample_completed_
      -- 
    ra_5498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2256_inst_ack_0, ack => convTransposeC_CP_4929_elements(60)); -- 
    -- CP-element group 61:  transition  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	57 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_1969/assign_stmt_2243_to_assign_stmt_2279/type_cast_2256_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_1969/assign_stmt_2243_to_assign_stmt_2279/type_cast_2256_Update/ca
      -- CP-element group 61: 	 branch_block_stmt_1969/assign_stmt_2243_to_assign_stmt_2279/type_cast_2273_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_1969/assign_stmt_2243_to_assign_stmt_2279/type_cast_2256_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_1969/assign_stmt_2243_to_assign_stmt_2279/type_cast_2273_Sample/rr
      -- CP-element group 61: 	 branch_block_stmt_1969/assign_stmt_2243_to_assign_stmt_2279/type_cast_2273_Sample/$entry
      -- 
    ca_5503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2256_inst_ack_1, ack => convTransposeC_CP_4929_elements(61)); -- 
    rr_5511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(61), ack => type_cast_2273_inst_req_0); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_1969/assign_stmt_2243_to_assign_stmt_2279/type_cast_2273_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_1969/assign_stmt_2243_to_assign_stmt_2279/type_cast_2273_Sample/ra
      -- CP-element group 62: 	 branch_block_stmt_1969/assign_stmt_2243_to_assign_stmt_2279/type_cast_2273_Sample/$exit
      -- 
    ra_5512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2273_inst_ack_0, ack => convTransposeC_CP_4929_elements(62)); -- 
    -- CP-element group 63:  branch  transition  place  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (13) 
      -- CP-element group 63: 	 branch_block_stmt_1969/assign_stmt_2243_to_assign_stmt_2279__exit__
      -- CP-element group 63: 	 branch_block_stmt_1969/assign_stmt_2243_to_assign_stmt_2279/type_cast_2273_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_1969/if_stmt_2280__entry__
      -- CP-element group 63: 	 branch_block_stmt_1969/assign_stmt_2243_to_assign_stmt_2279/type_cast_2273_Update/ca
      -- CP-element group 63: 	 branch_block_stmt_1969/if_stmt_2280_dead_link/$entry
      -- CP-element group 63: 	 branch_block_stmt_1969/if_stmt_2280_eval_test/$entry
      -- CP-element group 63: 	 branch_block_stmt_1969/assign_stmt_2243_to_assign_stmt_2279/$exit
      -- CP-element group 63: 	 branch_block_stmt_1969/if_stmt_2280_else_link/$entry
      -- CP-element group 63: 	 branch_block_stmt_1969/if_stmt_2280_if_link/$entry
      -- CP-element group 63: 	 branch_block_stmt_1969/R_cmp128_2281_place
      -- CP-element group 63: 	 branch_block_stmt_1969/assign_stmt_2243_to_assign_stmt_2279/type_cast_2273_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_1969/if_stmt_2280_eval_test/branch_req
      -- CP-element group 63: 	 branch_block_stmt_1969/if_stmt_2280_eval_test/$exit
      -- 
    ca_5517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2273_inst_ack_1, ack => convTransposeC_CP_4929_elements(63)); -- 
    branch_req_5525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(63), ack => if_stmt_2280_branch_req_0); -- 
    -- CP-element group 64:  merge  transition  place  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (15) 
      -- CP-element group 64: 	 branch_block_stmt_1969/merge_stmt_2286__exit__
      -- CP-element group 64: 	 branch_block_stmt_1969/assign_stmt_2291__entry__
      -- CP-element group 64: 	 branch_block_stmt_1969/merge_stmt_2286_PhiReqMerge
      -- CP-element group 64: 	 branch_block_stmt_1969/assign_stmt_2291/WPIPE_Block2_done_2288_Sample/req
      -- CP-element group 64: 	 branch_block_stmt_1969/assign_stmt_2291/WPIPE_Block2_done_2288_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_1969/assign_stmt_2291/WPIPE_Block2_done_2288_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_1969/assign_stmt_2291/$entry
      -- CP-element group 64: 	 branch_block_stmt_1969/ifx_xelse_whilex_xend
      -- CP-element group 64: 	 branch_block_stmt_1969/if_stmt_2280_if_link/if_choice_transition
      -- CP-element group 64: 	 branch_block_stmt_1969/if_stmt_2280_if_link/$exit
      -- CP-element group 64: 	 branch_block_stmt_1969/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 64: 	 branch_block_stmt_1969/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 64: 	 branch_block_stmt_1969/merge_stmt_2286_PhiAck/$entry
      -- CP-element group 64: 	 branch_block_stmt_1969/merge_stmt_2286_PhiAck/$exit
      -- CP-element group 64: 	 branch_block_stmt_1969/merge_stmt_2286_PhiAck/dummy
      -- 
    if_choice_transition_5530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2280_branch_ack_1, ack => convTransposeC_CP_4929_elements(64)); -- 
    req_5547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(64), ack => WPIPE_Block2_done_2288_inst_req_0); -- 
    -- CP-element group 65:  fork  transition  place  input  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	73 
    -- CP-element group 65: 	74 
    -- CP-element group 65: 	76 
    -- CP-element group 65: 	77 
    -- CP-element group 65:  members (20) 
      -- CP-element group 65: 	 branch_block_stmt_1969/ifx_xelse_whilex_xbodyx_xouter
      -- CP-element group 65: 	 branch_block_stmt_1969/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/type_cast_2061/SplitProtocol/Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1969/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/type_cast_2067/SplitProtocol/Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_1969/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/type_cast_2067/SplitProtocol/Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1969/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 65: 	 branch_block_stmt_1969/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/type_cast_2061/$entry
      -- CP-element group 65: 	 branch_block_stmt_1969/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2062/$entry
      -- CP-element group 65: 	 branch_block_stmt_1969/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/type_cast_2061/SplitProtocol/Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1969/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/$entry
      -- CP-element group 65: 	 branch_block_stmt_1969/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/type_cast_2067/$entry
      -- CP-element group 65: 	 branch_block_stmt_1969/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2055/$entry
      -- CP-element group 65: 	 branch_block_stmt_1969/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/type_cast_2067/SplitProtocol/$entry
      -- CP-element group 65: 	 branch_block_stmt_1969/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/type_cast_2067/SplitProtocol/Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1969/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/type_cast_2061/SplitProtocol/Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_1969/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/type_cast_2061/SplitProtocol/Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_1969/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/type_cast_2061/SplitProtocol/$entry
      -- CP-element group 65: 	 branch_block_stmt_1969/if_stmt_2280_else_link/else_choice_transition
      -- CP-element group 65: 	 branch_block_stmt_1969/if_stmt_2280_else_link/$exit
      -- CP-element group 65: 	 branch_block_stmt_1969/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/$entry
      -- CP-element group 65: 	 branch_block_stmt_1969/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/type_cast_2067/SplitProtocol/Sample/$entry
      -- 
    else_choice_transition_5534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2280_branch_ack_0, ack => convTransposeC_CP_4929_elements(65)); -- 
    rr_5606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(65), ack => type_cast_2067_inst_req_0); -- 
    cr_5634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(65), ack => type_cast_2061_inst_req_1); -- 
    cr_5611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(65), ack => type_cast_2067_inst_req_1); -- 
    rr_5629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(65), ack => type_cast_2061_inst_req_0); -- 
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_1969/assign_stmt_2291/WPIPE_Block2_done_2288_Update/req
      -- CP-element group 66: 	 branch_block_stmt_1969/assign_stmt_2291/WPIPE_Block2_done_2288_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_1969/assign_stmt_2291/WPIPE_Block2_done_2288_Sample/ack
      -- CP-element group 66: 	 branch_block_stmt_1969/assign_stmt_2291/WPIPE_Block2_done_2288_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_1969/assign_stmt_2291/WPIPE_Block2_done_2288_update_start_
      -- CP-element group 66: 	 branch_block_stmt_1969/assign_stmt_2291/WPIPE_Block2_done_2288_sample_completed_
      -- 
    ack_5548_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2288_inst_ack_0, ack => convTransposeC_CP_4929_elements(66)); -- 
    req_5552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(66), ack => WPIPE_Block2_done_2288_inst_req_1); -- 
    -- CP-element group 67:  transition  place  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (16) 
      -- CP-element group 67: 	 branch_block_stmt_1969/return__
      -- CP-element group 67: 	 branch_block_stmt_1969/assign_stmt_2291__exit__
      -- CP-element group 67: 	 $exit
      -- CP-element group 67: 	 branch_block_stmt_1969/$exit
      -- CP-element group 67: 	 branch_block_stmt_1969/merge_stmt_2293__exit__
      -- CP-element group 67: 	 branch_block_stmt_1969/branch_block_stmt_1969__exit__
      -- CP-element group 67: 	 branch_block_stmt_1969/merge_stmt_2293_PhiReqMerge
      -- CP-element group 67: 	 branch_block_stmt_1969/assign_stmt_2291/WPIPE_Block2_done_2288_Update/ack
      -- CP-element group 67: 	 branch_block_stmt_1969/assign_stmt_2291/WPIPE_Block2_done_2288_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_1969/assign_stmt_2291/WPIPE_Block2_done_2288_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_1969/assign_stmt_2291/$exit
      -- CP-element group 67: 	 branch_block_stmt_1969/return___PhiReq/$entry
      -- CP-element group 67: 	 branch_block_stmt_1969/return___PhiReq/$exit
      -- CP-element group 67: 	 branch_block_stmt_1969/merge_stmt_2293_PhiAck/$entry
      -- CP-element group 67: 	 branch_block_stmt_1969/merge_stmt_2293_PhiAck/$exit
      -- CP-element group 67: 	 branch_block_stmt_1969/merge_stmt_2293_PhiAck/dummy
      -- 
    ack_5553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2288_inst_ack_1, ack => convTransposeC_CP_4929_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	31 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (2) 
      -- CP-element group 68: 	 branch_block_stmt_1969/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/type_cast_2065/SplitProtocol/Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_1969/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/type_cast_2065/SplitProtocol/Sample/ra
      -- 
    ra_5573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2065_inst_ack_0, ack => convTransposeC_CP_4929_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	31 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (2) 
      -- CP-element group 69: 	 branch_block_stmt_1969/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/type_cast_2065/SplitProtocol/Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_1969/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/type_cast_2065/SplitProtocol/Update/ca
      -- 
    ca_5578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2065_inst_ack_1, ack => convTransposeC_CP_4929_elements(69)); -- 
    -- CP-element group 70:  join  transition  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (5) 
      -- CP-element group 70: 	 branch_block_stmt_1969/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/type_cast_2065/$exit
      -- CP-element group 70: 	 branch_block_stmt_1969/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/type_cast_2065/SplitProtocol/$exit
      -- CP-element group 70: 	 branch_block_stmt_1969/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2062/phi_stmt_2062_req
      -- CP-element group 70: 	 branch_block_stmt_1969/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/$exit
      -- CP-element group 70: 	 branch_block_stmt_1969/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2062/$exit
      -- 
    phi_stmt_2062_req_5579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2062_req_5579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(70), ack => phi_stmt_2062_req_0); -- 
    convTransposeC_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_4929_elements(68) & convTransposeC_CP_4929_elements(69);
      gj_convTransposeC_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_4929_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  transition  output  delay-element  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	31 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (4) 
      -- CP-element group 71: 	 branch_block_stmt_1969/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2055/$exit
      -- CP-element group 71: 	 branch_block_stmt_1969/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/$exit
      -- CP-element group 71: 	 branch_block_stmt_1969/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/type_cast_2059_konst_delay_trans
      -- CP-element group 71: 	 branch_block_stmt_1969/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2055/phi_stmt_2055_req
      -- 
    phi_stmt_2055_req_5587_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2055_req_5587_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(71), ack => phi_stmt_2055_req_0); -- 
    -- Element group convTransposeC_CP_4929_elements(71) is a control-delay.
    cp_element_71_delay: control_delay_element  generic map(name => " 71_delay", delay_value => 1)  port map(req => convTransposeC_CP_4929_elements(31), ack => convTransposeC_CP_4929_elements(71), clk => clk, reset =>reset);
    -- CP-element group 72:  join  transition  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	80 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_1969/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_4929_elements(70) & convTransposeC_CP_4929_elements(71);
      gj_convTransposeC_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_4929_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	65 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (2) 
      -- CP-element group 73: 	 branch_block_stmt_1969/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/type_cast_2067/SplitProtocol/Sample/ra
      -- CP-element group 73: 	 branch_block_stmt_1969/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/type_cast_2067/SplitProtocol/Sample/$exit
      -- 
    ra_5607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2067_inst_ack_0, ack => convTransposeC_CP_4929_elements(73)); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	65 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74:  members (2) 
      -- CP-element group 74: 	 branch_block_stmt_1969/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/type_cast_2067/SplitProtocol/Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_1969/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/type_cast_2067/SplitProtocol/Update/ca
      -- 
    ca_5612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2067_inst_ack_1, ack => convTransposeC_CP_4929_elements(74)); -- 
    -- CP-element group 75:  join  transition  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	79 
    -- CP-element group 75:  members (5) 
      -- CP-element group 75: 	 branch_block_stmt_1969/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2062/phi_stmt_2062_req
      -- CP-element group 75: 	 branch_block_stmt_1969/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2062/$exit
      -- CP-element group 75: 	 branch_block_stmt_1969/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/$exit
      -- CP-element group 75: 	 branch_block_stmt_1969/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/type_cast_2067/$exit
      -- CP-element group 75: 	 branch_block_stmt_1969/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2062/phi_stmt_2062_sources/type_cast_2067/SplitProtocol/$exit
      -- 
    phi_stmt_2062_req_5613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2062_req_5613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(75), ack => phi_stmt_2062_req_1); -- 
    convTransposeC_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_4929_elements(73) & convTransposeC_CP_4929_elements(74);
      gj_convTransposeC_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_4929_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	65 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (2) 
      -- CP-element group 76: 	 branch_block_stmt_1969/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/type_cast_2061/SplitProtocol/Sample/ra
      -- CP-element group 76: 	 branch_block_stmt_1969/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/type_cast_2061/SplitProtocol/Sample/$exit
      -- 
    ra_5630_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2061_inst_ack_0, ack => convTransposeC_CP_4929_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	65 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_1969/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/type_cast_2061/SplitProtocol/Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_1969/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/type_cast_2061/SplitProtocol/Update/ca
      -- 
    ca_5635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2061_inst_ack_1, ack => convTransposeC_CP_4929_elements(77)); -- 
    -- CP-element group 78:  join  transition  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (5) 
      -- CP-element group 78: 	 branch_block_stmt_1969/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2055/$exit
      -- CP-element group 78: 	 branch_block_stmt_1969/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2055/phi_stmt_2055_req
      -- CP-element group 78: 	 branch_block_stmt_1969/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/$exit
      -- CP-element group 78: 	 branch_block_stmt_1969/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/type_cast_2061/SplitProtocol/$exit
      -- CP-element group 78: 	 branch_block_stmt_1969/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/type_cast_2061/$exit
      -- 
    phi_stmt_2055_req_5636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2055_req_5636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(78), ack => phi_stmt_2055_req_1); -- 
    convTransposeC_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_4929_elements(76) & convTransposeC_CP_4929_elements(77);
      gj_convTransposeC_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_4929_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  join  transition  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	75 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_1969/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_4929_elements(75) & convTransposeC_CP_4929_elements(78);
      gj_convTransposeC_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_4929_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  merge  fork  transition  place  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	72 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_1969/merge_stmt_2054_PhiReqMerge
      -- CP-element group 80: 	 branch_block_stmt_1969/merge_stmt_2054_PhiAck/$entry
      -- 
    convTransposeC_CP_4929_elements(80) <= OrReduce(convTransposeC_CP_4929_elements(72) & convTransposeC_CP_4929_elements(79));
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_1969/merge_stmt_2054_PhiAck/phi_stmt_2055_ack
      -- 
    phi_stmt_2055_ack_5641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2055_ack_0, ack => convTransposeC_CP_4929_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_1969/merge_stmt_2054_PhiAck/phi_stmt_2062_ack
      -- 
    phi_stmt_2062_ack_5642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2062_ack_0, ack => convTransposeC_CP_4929_elements(82)); -- 
    -- CP-element group 83:  join  transition  place  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	87 
    -- CP-element group 83:  members (10) 
      -- CP-element group 83: 	 branch_block_stmt_1969/assign_stmt_2073_to_assign_stmt_2118__exit__
      -- CP-element group 83: 	 branch_block_stmt_1969/merge_stmt_2054__exit__
      -- CP-element group 83: 	 branch_block_stmt_1969/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 83: 	 branch_block_stmt_1969/assign_stmt_2073_to_assign_stmt_2118__entry__
      -- CP-element group 83: 	 branch_block_stmt_1969/merge_stmt_2054_PhiAck/$exit
      -- CP-element group 83: 	 branch_block_stmt_1969/assign_stmt_2073_to_assign_stmt_2118/$entry
      -- CP-element group 83: 	 branch_block_stmt_1969/assign_stmt_2073_to_assign_stmt_2118/$exit
      -- CP-element group 83: 	 branch_block_stmt_1969/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- CP-element group 83: 	 branch_block_stmt_1969/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2121/$entry
      -- CP-element group 83: 	 branch_block_stmt_1969/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2121/phi_stmt_2121_sources/$entry
      -- 
    convTransposeC_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_4929_elements(81) & convTransposeC_CP_4929_elements(82);
      gj_convTransposeC_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_4929_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	56 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_1969/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2121/phi_stmt_2121_sources/type_cast_2127/SplitProtocol/Sample/ra
      -- CP-element group 84: 	 branch_block_stmt_1969/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2121/phi_stmt_2121_sources/type_cast_2127/SplitProtocol/Sample/$exit
      -- 
    ra_5662_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2127_inst_ack_0, ack => convTransposeC_CP_4929_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	56 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_1969/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2121/phi_stmt_2121_sources/type_cast_2127/SplitProtocol/Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_1969/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2121/phi_stmt_2121_sources/type_cast_2127/SplitProtocol/Update/ca
      -- 
    ca_5667_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2127_inst_ack_1, ack => convTransposeC_CP_4929_elements(85)); -- 
    -- CP-element group 86:  join  transition  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (6) 
      -- CP-element group 86: 	 branch_block_stmt_1969/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2121/$exit
      -- CP-element group 86: 	 branch_block_stmt_1969/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2121/phi_stmt_2121_sources/$exit
      -- CP-element group 86: 	 branch_block_stmt_1969/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2121/phi_stmt_2121_sources/type_cast_2127/SplitProtocol/$exit
      -- CP-element group 86: 	 branch_block_stmt_1969/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2121/phi_stmt_2121_sources/type_cast_2127/$exit
      -- CP-element group 86: 	 branch_block_stmt_1969/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- CP-element group 86: 	 branch_block_stmt_1969/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2121/phi_stmt_2121_req
      -- 
    phi_stmt_2121_req_5668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2121_req_5668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(86), ack => phi_stmt_2121_req_1); -- 
    convTransposeC_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_4929_elements(84) & convTransposeC_CP_4929_elements(85);
      gj_convTransposeC_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_4929_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  transition  output  delay-element  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	83 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (5) 
      -- CP-element group 87: 	 branch_block_stmt_1969/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- CP-element group 87: 	 branch_block_stmt_1969/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2121/$exit
      -- CP-element group 87: 	 branch_block_stmt_1969/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2121/phi_stmt_2121_sources/$exit
      -- CP-element group 87: 	 branch_block_stmt_1969/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2121/phi_stmt_2121_sources/type_cast_2125_konst_delay_trans
      -- CP-element group 87: 	 branch_block_stmt_1969/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2121/phi_stmt_2121_req
      -- 
    phi_stmt_2121_req_5679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2121_req_5679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(87), ack => phi_stmt_2121_req_0); -- 
    -- Element group convTransposeC_CP_4929_elements(87) is a control-delay.
    cp_element_87_delay: control_delay_element  generic map(name => " 87_delay", delay_value => 1)  port map(req => convTransposeC_CP_4929_elements(83), ack => convTransposeC_CP_4929_elements(87), clk => clk, reset =>reset);
    -- CP-element group 88:  merge  transition  place  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_1969/merge_stmt_2120_PhiReqMerge
      -- CP-element group 88: 	 branch_block_stmt_1969/merge_stmt_2120_PhiAck/$entry
      -- 
    convTransposeC_CP_4929_elements(88) <= OrReduce(convTransposeC_CP_4929_elements(86) & convTransposeC_CP_4929_elements(87));
    -- CP-element group 89:  fork  transition  place  input  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	32 
    -- CP-element group 89: 	33 
    -- CP-element group 89: 	35 
    -- CP-element group 89: 	37 
    -- CP-element group 89: 	39 
    -- CP-element group 89: 	41 
    -- CP-element group 89: 	42 
    -- CP-element group 89: 	43 
    -- CP-element group 89: 	45 
    -- CP-element group 89: 	47 
    -- CP-element group 89: 	49 
    -- CP-element group 89: 	52 
    -- CP-element group 89: 	53 
    -- CP-element group 89: 	54 
    -- CP-element group 89:  members (51) 
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2168_final_index_sum_regn_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222__entry__
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2168_final_index_sum_regn_Update/req
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2178_Update/cr
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2198_final_index_sum_regn_update_start
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2173_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2208_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_1969/merge_stmt_2120__exit__
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2208_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2202_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2208_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2198_final_index_sum_regn_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2173_Update/word_access_complete/$entry
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2208_Sample/rr
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2173_Update/word_access_complete/word_0/$entry
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2173_Update/word_access_complete/word_0/cr
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2198_final_index_sum_regn_Update/req
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2178_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2208_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2192_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2208_Update/cr
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2178_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2178_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2178_Sample/rr
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/addr_of_2199_complete/$entry
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/addr_of_2199_complete/req
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/addr_of_2169_complete/$entry
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2202_Update/word_access_complete/word_0/cr
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2173_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2202_Update/word_access_complete/word_0/$entry
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2202_Update/word_access_complete/$entry
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/ptr_deref_2202_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/addr_of_2199_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/addr_of_2169_complete/req
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2192_Update/cr
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2192_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/$entry
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2148_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2148_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2148_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2178_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2148_Sample/rr
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2148_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2148_Update/cr
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2162_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2162_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/type_cast_2162_Update/cr
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/addr_of_2169_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1969/assign_stmt_2134_to_assign_stmt_2222/array_obj_ref_2168_final_index_sum_regn_update_start
      -- CP-element group 89: 	 branch_block_stmt_1969/merge_stmt_2120_PhiAck/$exit
      -- CP-element group 89: 	 branch_block_stmt_1969/merge_stmt_2120_PhiAck/phi_stmt_2121_ack
      -- 
    phi_stmt_2121_ack_5684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2121_ack_0, ack => convTransposeC_CP_4929_elements(89)); -- 
    req_5246_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5246_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(89), ack => array_obj_ref_2168_index_offset_req_1); -- 
    cr_5325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(89), ack => type_cast_2178_inst_req_1); -- 
    rr_5444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(89), ack => type_cast_2208_inst_req_0); -- 
    cr_5306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(89), ack => ptr_deref_2173_load_0_req_1); -- 
    req_5370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(89), ack => array_obj_ref_2198_index_offset_req_1); -- 
    cr_5449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(89), ack => type_cast_2208_inst_req_1); -- 
    rr_5320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(89), ack => type_cast_2178_inst_req_0); -- 
    req_5385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(89), ack => addr_of_2199_final_reg_req_1); -- 
    cr_5435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(89), ack => ptr_deref_2202_store_0_req_1); -- 
    req_5261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(89), ack => addr_of_2169_final_reg_req_1); -- 
    cr_5339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(89), ack => type_cast_2192_inst_req_1); -- 
    rr_5196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(89), ack => type_cast_2148_inst_req_0); -- 
    cr_5201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(89), ack => type_cast_2148_inst_req_1); -- 
    cr_5215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4929_elements(89), ack => type_cast_2162_inst_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_2156_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2186_wire : std_logic_vector(31 downto 0);
    signal R_idxprom97_2197_resized : std_logic_vector(13 downto 0);
    signal R_idxprom97_2197_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2167_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2167_scaled : std_logic_vector(13 downto 0);
    signal add102_2215 : std_logic_vector(31 downto 0);
    signal add44_2139 : std_logic_vector(15 downto 0);
    signal add88_2144 : std_logic_vector(15 downto 0);
    signal array_obj_ref_2168_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2168_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2168_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2168_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2168_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2168_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2198_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2198_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2198_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2198_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2198_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2198_root_address : std_logic_vector(13 downto 0);
    signal arrayidx92_2170 : std_logic_vector(31 downto 0);
    signal arrayidx98_2200 : std_logic_vector(31 downto 0);
    signal call11_1990 : std_logic_vector(15 downto 0);
    signal call13_1993 : std_logic_vector(15 downto 0);
    signal call14_1996 : std_logic_vector(15 downto 0);
    signal call15_1999 : std_logic_vector(15 downto 0);
    signal call17_2002 : std_logic_vector(15 downto 0);
    signal call19_2005 : std_logic_vector(15 downto 0);
    signal call1_1975 : std_logic_vector(15 downto 0);
    signal call3_1978 : std_logic_vector(15 downto 0);
    signal call5_1981 : std_logic_vector(15 downto 0);
    signal call7_1984 : std_logic_vector(15 downto 0);
    signal call9_1987 : std_logic_vector(15 downto 0);
    signal call_1972 : std_logic_vector(15 downto 0);
    signal cmp118_2253 : std_logic_vector(0 downto 0);
    signal cmp128_2279 : std_logic_vector(0 downto 0);
    signal cmp_2222 : std_logic_vector(0 downto 0);
    signal conv101_2209 : std_logic_vector(31 downto 0);
    signal conv105_2016 : std_logic_vector(31 downto 0);
    signal conv113_2248 : std_logic_vector(31 downto 0);
    signal conv116_2020 : std_logic_vector(31 downto 0);
    signal conv124_2274 : std_logic_vector(31 downto 0);
    signal conv127_2030 : std_logic_vector(31 downto 0);
    signal conv91_2149 : std_logic_vector(31 downto 0);
    signal conv95_2179 : std_logic_vector(31 downto 0);
    signal div117_2026 : std_logic_vector(31 downto 0);
    signal div_2012 : std_logic_vector(15 downto 0);
    signal idxprom97_2193 : std_logic_vector(63 downto 0);
    signal idxprom_2163 : std_logic_vector(63 downto 0);
    signal inc122_2257 : std_logic_vector(15 downto 0);
    signal inc122x_xinput_dim0x_x2_2262 : std_logic_vector(15 downto 0);
    signal inc_2243 : std_logic_vector(15 downto 0);
    signal indvar_2121 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_2235 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_2062 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_2055 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2269 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2134 : std_logic_vector(15 downto 0);
    signal ptr_deref_2173_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2173_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2173_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2173_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2173_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2202_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2202_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2202_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2202_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2202_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2202_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr96_2188 : std_logic_vector(31 downto 0);
    signal shr_2158 : std_logic_vector(31 downto 0);
    signal tmp10_2118 : std_logic_vector(15 downto 0);
    signal tmp155_2073 : std_logic_vector(15 downto 0);
    signal tmp156_2078 : std_logic_vector(15 downto 0);
    signal tmp157_2083 : std_logic_vector(15 downto 0);
    signal tmp1_2041 : std_logic_vector(15 downto 0);
    signal tmp2_2088 : std_logic_vector(15 downto 0);
    signal tmp3_2093 : std_logic_vector(15 downto 0);
    signal tmp4_2047 : std_logic_vector(15 downto 0);
    signal tmp5_2052 : std_logic_vector(15 downto 0);
    signal tmp6_2098 : std_logic_vector(15 downto 0);
    signal tmp7_2103 : std_logic_vector(15 downto 0);
    signal tmp8_2108 : std_logic_vector(15 downto 0);
    signal tmp93_2174 : std_logic_vector(63 downto 0);
    signal tmp9_2113 : std_logic_vector(15 downto 0);
    signal tmp_2036 : std_logic_vector(15 downto 0);
    signal type_cast_2010_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2024_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2034_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2045_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2059_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2061_wire : std_logic_vector(15 downto 0);
    signal type_cast_2065_wire : std_logic_vector(15 downto 0);
    signal type_cast_2067_wire : std_logic_vector(15 downto 0);
    signal type_cast_2125_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2127_wire : std_logic_vector(15 downto 0);
    signal type_cast_2132_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2147_wire : std_logic_vector(31 downto 0);
    signal type_cast_2152_wire : std_logic_vector(31 downto 0);
    signal type_cast_2155_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2161_wire : std_logic_vector(63 downto 0);
    signal type_cast_2177_wire : std_logic_vector(31 downto 0);
    signal type_cast_2182_wire : std_logic_vector(31 downto 0);
    signal type_cast_2185_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2191_wire : std_logic_vector(63 downto 0);
    signal type_cast_2207_wire : std_logic_vector(31 downto 0);
    signal type_cast_2213_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2218_wire : std_logic_vector(31 downto 0);
    signal type_cast_2220_wire : std_logic_vector(31 downto 0);
    signal type_cast_2233_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2241_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2246_wire : std_logic_vector(31 downto 0);
    signal type_cast_2266_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2272_wire : std_logic_vector(31 downto 0);
    signal type_cast_2290_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_2168_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2168_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2168_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2168_resized_base_address <= "00000000000000";
    array_obj_ref_2198_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2198_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2198_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2198_resized_base_address <= "00000000000000";
    ptr_deref_2173_word_offset_0 <= "00000000000000";
    ptr_deref_2202_word_offset_0 <= "00000000000000";
    type_cast_2010_wire_constant <= "0000000000000001";
    type_cast_2024_wire_constant <= "00000000000000000000000000000001";
    type_cast_2034_wire_constant <= "1111111111111111";
    type_cast_2045_wire_constant <= "1111111111111111";
    type_cast_2059_wire_constant <= "0000000000000000";
    type_cast_2125_wire_constant <= "0000000000000000";
    type_cast_2132_wire_constant <= "0000000000000100";
    type_cast_2155_wire_constant <= "00000000000000000000000000000010";
    type_cast_2185_wire_constant <= "00000000000000000000000000000010";
    type_cast_2213_wire_constant <= "00000000000000000000000000000100";
    type_cast_2233_wire_constant <= "0000000000000001";
    type_cast_2241_wire_constant <= "0000000000000001";
    type_cast_2266_wire_constant <= "0000000000000000";
    type_cast_2290_wire_constant <= "0000000000000001";
    phi_stmt_2055: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2059_wire_constant & type_cast_2061_wire;
      req <= phi_stmt_2055_req_0 & phi_stmt_2055_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2055",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2055_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_2055,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2055
    phi_stmt_2062: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2065_wire & type_cast_2067_wire;
      req <= phi_stmt_2062_req_0 & phi_stmt_2062_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2062",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2062_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_2062,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2062
    phi_stmt_2121: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2125_wire_constant & type_cast_2127_wire;
      req <= phi_stmt_2121_req_0 & phi_stmt_2121_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2121",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2121_ack_0,
          idata => idata,
          odata => indvar_2121,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2121
    -- flow-through select operator MUX_2268_inst
    input_dim1x_x2_2269 <= type_cast_2266_wire_constant when (cmp118_2253(0) /=  '0') else inc_2243;
    addr_of_2169_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2169_final_reg_req_0;
      addr_of_2169_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2169_final_reg_req_1;
      addr_of_2169_final_reg_ack_1<= rack(0);
      addr_of_2169_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2169_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2168_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx92_2170,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2199_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2199_final_reg_req_0;
      addr_of_2199_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2199_final_reg_req_1;
      addr_of_2199_final_reg_ack_1<= rack(0);
      addr_of_2199_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2199_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2198_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx98_2200,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2015_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2015_inst_req_0;
      type_cast_2015_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2015_inst_req_1;
      type_cast_2015_inst_ack_1<= rack(0);
      type_cast_2015_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2015_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_1978,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv105_2016,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2019_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2019_inst_req_0;
      type_cast_2019_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2019_inst_req_1;
      type_cast_2019_inst_ack_1<= rack(0);
      type_cast_2019_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2019_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1_1975,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv116_2020,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2029_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2029_inst_req_0;
      type_cast_2029_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2029_inst_req_1;
      type_cast_2029_inst_ack_1<= rack(0);
      type_cast_2029_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2029_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1972,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv127_2030,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2061_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2061_inst_req_0;
      type_cast_2061_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2061_inst_req_1;
      type_cast_2061_inst_ack_1<= rack(0);
      type_cast_2061_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2061_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2269,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2061_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2065_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2065_inst_req_0;
      type_cast_2065_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2065_inst_req_1;
      type_cast_2065_inst_ack_1<= rack(0);
      type_cast_2065_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2065_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_2012,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2065_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2067_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2067_inst_req_0;
      type_cast_2067_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2067_inst_req_1;
      type_cast_2067_inst_ack_1<= rack(0);
      type_cast_2067_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2067_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc122x_xinput_dim0x_x2_2262,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2067_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2127_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2127_inst_req_0;
      type_cast_2127_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2127_inst_req_1;
      type_cast_2127_inst_ack_1<= rack(0);
      type_cast_2127_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2127_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2235,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2127_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2148_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2148_inst_req_0;
      type_cast_2148_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2148_inst_req_1;
      type_cast_2148_inst_ack_1<= rack(0);
      type_cast_2148_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2148_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2147_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv91_2149,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2152_inst
    process(conv91_2149) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv91_2149(31 downto 0);
      type_cast_2152_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2157_inst
    process(ASHR_i32_i32_2156_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2156_wire(31 downto 0);
      shr_2158 <= tmp_var; -- 
    end process;
    type_cast_2162_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2162_inst_req_0;
      type_cast_2162_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2162_inst_req_1;
      type_cast_2162_inst_ack_1<= rack(0);
      type_cast_2162_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2162_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2161_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2163,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2178_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2178_inst_req_0;
      type_cast_2178_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2178_inst_req_1;
      type_cast_2178_inst_ack_1<= rack(0);
      type_cast_2178_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2178_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2177_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_2179,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2182_inst
    process(conv95_2179) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv95_2179(31 downto 0);
      type_cast_2182_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2187_inst
    process(ASHR_i32_i32_2186_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2186_wire(31 downto 0);
      shr96_2188 <= tmp_var; -- 
    end process;
    type_cast_2192_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2192_inst_req_0;
      type_cast_2192_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2192_inst_req_1;
      type_cast_2192_inst_ack_1<= rack(0);
      type_cast_2192_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2192_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2191_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom97_2193,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2208_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2208_inst_req_0;
      type_cast_2208_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2208_inst_req_1;
      type_cast_2208_inst_ack_1<= rack(0);
      type_cast_2208_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2208_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2207_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv101_2209,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2218_inst
    process(add102_2215) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add102_2215(31 downto 0);
      type_cast_2218_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2220_inst
    process(conv105_2016) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv105_2016(31 downto 0);
      type_cast_2220_wire <= tmp_var; -- 
    end process;
    type_cast_2247_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2247_inst_req_0;
      type_cast_2247_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2247_inst_req_1;
      type_cast_2247_inst_ack_1<= rack(0);
      type_cast_2247_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2247_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2246_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv113_2248,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2256_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2256_inst_req_0;
      type_cast_2256_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2256_inst_req_1;
      type_cast_2256_inst_ack_1<= rack(0);
      type_cast_2256_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2256_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp118_2253,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc122_2257,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2273_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2273_inst_req_0;
      type_cast_2273_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2273_inst_req_1;
      type_cast_2273_inst_ack_1<= rack(0);
      type_cast_2273_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2273_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2272_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv124_2274,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_2168_index_1_rename
    process(R_idxprom_2167_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2167_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2167_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2168_index_1_resize
    process(idxprom_2163) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2163;
      ov := iv(13 downto 0);
      R_idxprom_2167_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2168_root_address_inst
    process(array_obj_ref_2168_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2168_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2168_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2198_index_1_rename
    process(R_idxprom97_2197_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom97_2197_resized;
      ov(13 downto 0) := iv;
      R_idxprom97_2197_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2198_index_1_resize
    process(idxprom97_2193) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom97_2193;
      ov := iv(13 downto 0);
      R_idxprom97_2197_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2198_root_address_inst
    process(array_obj_ref_2198_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2198_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2198_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2173_addr_0
    process(ptr_deref_2173_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2173_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2173_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2173_base_resize
    process(arrayidx92_2170) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx92_2170;
      ov := iv(13 downto 0);
      ptr_deref_2173_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2173_gather_scatter
    process(ptr_deref_2173_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2173_data_0;
      ov(63 downto 0) := iv;
      tmp93_2174 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2173_root_address_inst
    process(ptr_deref_2173_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2173_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2173_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2202_addr_0
    process(ptr_deref_2202_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2202_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2202_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2202_base_resize
    process(arrayidx98_2200) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx98_2200;
      ov := iv(13 downto 0);
      ptr_deref_2202_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2202_gather_scatter
    process(tmp93_2174) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp93_2174;
      ov(63 downto 0) := iv;
      ptr_deref_2202_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2202_root_address_inst
    process(ptr_deref_2202_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2202_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2202_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2223_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2222;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2223_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2223_branch_req_0,
          ack0 => if_stmt_2223_branch_ack_0,
          ack1 => if_stmt_2223_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2280_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp128_2279;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2280_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2280_branch_req_0,
          ack0 => if_stmt_2280_branch_ack_0,
          ack1 => if_stmt_2280_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2035_inst
    process(call9_1987) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_1987, type_cast_2034_wire_constant, tmp_var);
      tmp_2036 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2046_inst
    process(call7_1984) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_1984, type_cast_2045_wire_constant, tmp_var);
      tmp4_2047 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2077_inst
    process(input_dim1x_x1x_xph_2055, tmp155_2073) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_2055, tmp155_2073, tmp_var);
      tmp156_2078 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2092_inst
    process(tmp1_2041, tmp2_2088) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp1_2041, tmp2_2088, tmp_var);
      tmp3_2093 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2102_inst
    process(tmp5_2052, tmp6_2098) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp5_2052, tmp6_2098, tmp_var);
      tmp7_2103 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2112_inst
    process(tmp3_2093, tmp8_2108) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp3_2093, tmp8_2108, tmp_var);
      tmp9_2113 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2138_inst
    process(tmp157_2083, input_dim2x_x1_2134) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp157_2083, input_dim2x_x1_2134, tmp_var);
      add44_2139 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2143_inst
    process(tmp10_2118, input_dim2x_x1_2134) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp10_2118, input_dim2x_x1_2134, tmp_var);
      add88_2144 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2234_inst
    process(indvar_2121) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2121, type_cast_2233_wire_constant, tmp_var);
      indvarx_xnext_2235 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2242_inst
    process(input_dim1x_x1x_xph_2055) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_2055, type_cast_2241_wire_constant, tmp_var);
      inc_2243 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2261_inst
    process(inc122_2257, input_dim0x_x2x_xph_2062) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc122_2257, input_dim0x_x2x_xph_2062, tmp_var);
      inc122x_xinput_dim0x_x2_2262 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2214_inst
    process(conv101_2209) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv101_2209, type_cast_2213_wire_constant, tmp_var);
      add102_2215 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2156_inst
    process(type_cast_2152_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2152_wire, type_cast_2155_wire_constant, tmp_var);
      ASHR_i32_i32_2156_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2186_inst
    process(type_cast_2182_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2182_wire, type_cast_2185_wire_constant, tmp_var);
      ASHR_i32_i32_2186_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2252_inst
    process(conv113_2248, div117_2026) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv113_2248, div117_2026, tmp_var);
      cmp118_2253 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2278_inst
    process(conv124_2274, conv127_2030) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv124_2274, conv127_2030, tmp_var);
      cmp128_2279 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2011_inst
    process(call_1972) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_1972, type_cast_2010_wire_constant, tmp_var);
      div_2012 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2025_inst
    process(conv116_2020) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv116_2020, type_cast_2024_wire_constant, tmp_var);
      div117_2026 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2072_inst
    process(call1_1975, input_dim0x_x2x_xph_2062) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call1_1975, input_dim0x_x2x_xph_2062, tmp_var);
      tmp155_2073 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2082_inst
    process(call3_1978, tmp156_2078) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call3_1978, tmp156_2078, tmp_var);
      tmp157_2083 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2087_inst
    process(call13_1993, input_dim1x_x1x_xph_2055) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call13_1993, input_dim1x_x1x_xph_2055, tmp_var);
      tmp2_2088 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2097_inst
    process(call13_1993, input_dim0x_x2x_xph_2062) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call13_1993, input_dim0x_x2x_xph_2062, tmp_var);
      tmp6_2098 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2107_inst
    process(call17_2002, tmp7_2103) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call17_2002, tmp7_2103, tmp_var);
      tmp8_2108 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2117_inst
    process(call19_2005, tmp9_2113) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call19_2005, tmp9_2113, tmp_var);
      tmp10_2118 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2133_inst
    process(indvar_2121) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2121, type_cast_2132_wire_constant, tmp_var);
      input_dim2x_x1_2134 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2221_inst
    process(type_cast_2218_wire, type_cast_2220_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2218_wire, type_cast_2220_wire, tmp_var);
      cmp_2222 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2040_inst
    process(tmp_2036, call14_1996) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp_2036, call14_1996, tmp_var);
      tmp1_2041 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2051_inst
    process(tmp4_2047, call14_1996) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp4_2047, call14_1996, tmp_var);
      tmp5_2052 <= tmp_var; --
    end process;
    -- shared split operator group (28) : array_obj_ref_2168_index_offset 
    ApIntAdd_group_28: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2167_scaled;
      array_obj_ref_2168_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2168_index_offset_req_0;
      array_obj_ref_2168_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2168_index_offset_req_1;
      array_obj_ref_2168_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_28_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_28_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : array_obj_ref_2198_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom97_2197_scaled;
      array_obj_ref_2198_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2198_index_offset_req_0;
      array_obj_ref_2198_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2198_index_offset_req_1;
      array_obj_ref_2198_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- unary operator type_cast_2147_inst
    process(add44_2139) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", add44_2139, tmp_var);
      type_cast_2147_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2161_inst
    process(shr_2158) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_2158, tmp_var);
      type_cast_2161_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2177_inst
    process(add88_2144) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", add88_2144, tmp_var);
      type_cast_2177_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2191_inst
    process(shr96_2188) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr96_2188, tmp_var);
      type_cast_2191_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2207_inst
    process(input_dim2x_x1_2134) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim2x_x1_2134, tmp_var);
      type_cast_2207_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2246_inst
    process(inc_2243) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_2243, tmp_var);
      type_cast_2246_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2272_inst
    process(inc122x_xinput_dim0x_x2_2262) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc122x_xinput_dim0x_x2_2262, tmp_var);
      type_cast_2272_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_2173_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2173_load_0_req_0;
      ptr_deref_2173_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2173_load_0_req_1;
      ptr_deref_2173_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2173_word_address_0;
      ptr_deref_2173_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_2202_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2202_store_0_req_0;
      ptr_deref_2202_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2202_store_0_req_1;
      ptr_deref_2202_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2202_word_address_0;
      data_in <= ptr_deref_2202_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block1_start_1971_inst RPIPE_Block1_start_1974_inst RPIPE_Block1_start_1977_inst RPIPE_Block1_start_1980_inst RPIPE_Block1_start_1983_inst RPIPE_Block1_start_1986_inst RPIPE_Block1_start_1989_inst RPIPE_Block1_start_1992_inst RPIPE_Block1_start_1995_inst RPIPE_Block1_start_1998_inst RPIPE_Block1_start_2001_inst RPIPE_Block1_start_2004_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(191 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 11 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 11 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 11 downto 0);
      signal guard_vector : std_logic_vector( 11 downto 0);
      constant outBUFs : IntegerArray(11 downto 0) := (11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(11 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false);
      constant guardBuffering: IntegerArray(11 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2);
      -- 
    begin -- 
      reqL_unguarded(11) <= RPIPE_Block1_start_1971_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block1_start_1974_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block1_start_1977_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block1_start_1980_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block1_start_1983_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block1_start_1986_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block1_start_1989_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block1_start_1992_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block1_start_1995_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block1_start_1998_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block1_start_2001_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block1_start_2004_inst_req_0;
      RPIPE_Block1_start_1971_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block1_start_1974_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block1_start_1977_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block1_start_1980_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block1_start_1983_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block1_start_1986_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block1_start_1989_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block1_start_1992_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block1_start_1995_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block1_start_1998_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block1_start_2001_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block1_start_2004_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(11) <= RPIPE_Block1_start_1971_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block1_start_1974_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block1_start_1977_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block1_start_1980_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block1_start_1983_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block1_start_1986_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block1_start_1989_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block1_start_1992_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block1_start_1995_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block1_start_1998_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block1_start_2001_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block1_start_2004_inst_req_1;
      RPIPE_Block1_start_1971_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block1_start_1974_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block1_start_1977_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block1_start_1980_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block1_start_1983_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block1_start_1986_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block1_start_1989_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block1_start_1992_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block1_start_1995_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block1_start_1998_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block1_start_2001_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block1_start_2004_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      call_1972 <= data_out(191 downto 176);
      call1_1975 <= data_out(175 downto 160);
      call3_1978 <= data_out(159 downto 144);
      call5_1981 <= data_out(143 downto 128);
      call7_1984 <= data_out(127 downto 112);
      call9_1987 <= data_out(111 downto 96);
      call11_1990 <= data_out(95 downto 80);
      call13_1993 <= data_out(79 downto 64);
      call14_1996 <= data_out(63 downto 48);
      call15_1999 <= data_out(47 downto 32);
      call17_2002 <= data_out(31 downto 16);
      call19_2005 <= data_out(15 downto 0);
      Block1_start_read_0_gI: SplitGuardInterface generic map(name => "Block1_start_read_0_gI", nreqs => 12, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_start_read_0: InputPortRevised -- 
        generic map ( name => "Block1_start_read_0", data_width => 16,  num_reqs => 12,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_start_pipe_read_req(0),
          oack => Block1_start_pipe_read_ack(0),
          odata => Block1_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block2_done_2288_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block2_done_2288_inst_req_0;
      WPIPE_Block2_done_2288_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block2_done_2288_inst_req_1;
      WPIPE_Block2_done_2288_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2290_wire_constant;
      Block2_done_write_0_gI: SplitGuardInterface generic map(name => "Block2_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block2_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_done_pipe_write_req(0),
          oack => Block2_done_pipe_write_ack(0),
          odata => Block2_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeC_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeD is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeD;
architecture convTransposeD_arch of convTransposeD is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeD_CP_5725_start: Boolean;
  signal convTransposeD_CP_5725_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block1_start_2299_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2299_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2302_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2299_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2299_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2302_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2302_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2302_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2305_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2308_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2308_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2305_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2308_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2311_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2311_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2305_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2308_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2305_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2311_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2311_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2314_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2314_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2314_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2314_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2317_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2317_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2317_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2317_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2320_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2320_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2320_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2320_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2323_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2323_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2323_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2323_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2326_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2326_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2326_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2326_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2329_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2329_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2329_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2329_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2332_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2332_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2332_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2332_inst_ack_1 : boolean;
  signal type_cast_2349_inst_req_0 : boolean;
  signal type_cast_2349_inst_ack_0 : boolean;
  signal type_cast_2349_inst_req_1 : boolean;
  signal type_cast_2349_inst_ack_1 : boolean;
  signal type_cast_2353_inst_req_0 : boolean;
  signal type_cast_2353_inst_ack_0 : boolean;
  signal type_cast_2353_inst_req_1 : boolean;
  signal type_cast_2353_inst_ack_1 : boolean;
  signal type_cast_2357_inst_req_0 : boolean;
  signal type_cast_2357_inst_ack_0 : boolean;
  signal type_cast_2357_inst_req_1 : boolean;
  signal type_cast_2357_inst_ack_1 : boolean;
  signal type_cast_2475_inst_req_0 : boolean;
  signal type_cast_2475_inst_ack_0 : boolean;
  signal type_cast_2475_inst_req_1 : boolean;
  signal type_cast_2475_inst_ack_1 : boolean;
  signal type_cast_2489_inst_req_0 : boolean;
  signal type_cast_2489_inst_ack_0 : boolean;
  signal type_cast_2489_inst_req_1 : boolean;
  signal type_cast_2489_inst_ack_1 : boolean;
  signal array_obj_ref_2495_index_offset_req_0 : boolean;
  signal array_obj_ref_2495_index_offset_ack_0 : boolean;
  signal array_obj_ref_2495_index_offset_req_1 : boolean;
  signal array_obj_ref_2495_index_offset_ack_1 : boolean;
  signal addr_of_2496_final_reg_req_0 : boolean;
  signal addr_of_2496_final_reg_ack_0 : boolean;
  signal addr_of_2496_final_reg_req_1 : boolean;
  signal addr_of_2496_final_reg_ack_1 : boolean;
  signal ptr_deref_2500_load_0_req_0 : boolean;
  signal ptr_deref_2500_load_0_ack_0 : boolean;
  signal ptr_deref_2500_load_0_req_1 : boolean;
  signal ptr_deref_2500_load_0_ack_1 : boolean;
  signal type_cast_2505_inst_req_0 : boolean;
  signal type_cast_2505_inst_ack_0 : boolean;
  signal type_cast_2505_inst_req_1 : boolean;
  signal type_cast_2505_inst_ack_1 : boolean;
  signal type_cast_2519_inst_req_0 : boolean;
  signal type_cast_2519_inst_ack_0 : boolean;
  signal type_cast_2519_inst_req_1 : boolean;
  signal type_cast_2519_inst_ack_1 : boolean;
  signal array_obj_ref_2525_index_offset_req_0 : boolean;
  signal array_obj_ref_2525_index_offset_ack_0 : boolean;
  signal array_obj_ref_2525_index_offset_req_1 : boolean;
  signal array_obj_ref_2525_index_offset_ack_1 : boolean;
  signal addr_of_2526_final_reg_req_0 : boolean;
  signal addr_of_2526_final_reg_ack_0 : boolean;
  signal addr_of_2526_final_reg_req_1 : boolean;
  signal addr_of_2526_final_reg_ack_1 : boolean;
  signal ptr_deref_2529_store_0_req_0 : boolean;
  signal ptr_deref_2529_store_0_ack_0 : boolean;
  signal ptr_deref_2529_store_0_req_1 : boolean;
  signal ptr_deref_2529_store_0_ack_1 : boolean;
  signal type_cast_2535_inst_req_0 : boolean;
  signal type_cast_2535_inst_ack_0 : boolean;
  signal type_cast_2535_inst_req_1 : boolean;
  signal type_cast_2535_inst_ack_1 : boolean;
  signal if_stmt_2550_branch_req_0 : boolean;
  signal if_stmt_2550_branch_ack_1 : boolean;
  signal if_stmt_2550_branch_ack_0 : boolean;
  signal type_cast_2574_inst_req_0 : boolean;
  signal type_cast_2574_inst_ack_0 : boolean;
  signal type_cast_2574_inst_req_1 : boolean;
  signal type_cast_2574_inst_ack_1 : boolean;
  signal type_cast_2589_inst_req_0 : boolean;
  signal type_cast_2589_inst_ack_0 : boolean;
  signal type_cast_2589_inst_req_1 : boolean;
  signal type_cast_2589_inst_ack_1 : boolean;
  signal type_cast_2599_inst_req_0 : boolean;
  signal type_cast_2599_inst_ack_0 : boolean;
  signal type_cast_2599_inst_req_1 : boolean;
  signal type_cast_2599_inst_ack_1 : boolean;
  signal if_stmt_2606_branch_req_0 : boolean;
  signal if_stmt_2606_branch_ack_1 : boolean;
  signal if_stmt_2606_branch_ack_0 : boolean;
  signal WPIPE_Block3_done_2614_inst_req_0 : boolean;
  signal WPIPE_Block3_done_2614_inst_ack_0 : boolean;
  signal WPIPE_Block3_done_2614_inst_req_1 : boolean;
  signal WPIPE_Block3_done_2614_inst_ack_1 : boolean;
  signal type_cast_2386_inst_req_0 : boolean;
  signal type_cast_2386_inst_ack_0 : boolean;
  signal type_cast_2386_inst_req_1 : boolean;
  signal type_cast_2386_inst_ack_1 : boolean;
  signal phi_stmt_2383_req_0 : boolean;
  signal type_cast_2394_inst_req_0 : boolean;
  signal type_cast_2394_inst_ack_0 : boolean;
  signal type_cast_2394_inst_req_1 : boolean;
  signal type_cast_2394_inst_ack_1 : boolean;
  signal phi_stmt_2389_req_1 : boolean;
  signal type_cast_2388_inst_req_0 : boolean;
  signal type_cast_2388_inst_ack_0 : boolean;
  signal type_cast_2388_inst_req_1 : boolean;
  signal type_cast_2388_inst_ack_1 : boolean;
  signal phi_stmt_2383_req_1 : boolean;
  signal type_cast_2392_inst_req_0 : boolean;
  signal type_cast_2392_inst_ack_0 : boolean;
  signal type_cast_2392_inst_req_1 : boolean;
  signal type_cast_2392_inst_ack_1 : boolean;
  signal phi_stmt_2389_req_0 : boolean;
  signal phi_stmt_2383_ack_0 : boolean;
  signal phi_stmt_2389_ack_0 : boolean;
  signal type_cast_2451_inst_req_0 : boolean;
  signal type_cast_2451_inst_ack_0 : boolean;
  signal type_cast_2451_inst_req_1 : boolean;
  signal type_cast_2451_inst_ack_1 : boolean;
  signal phi_stmt_2448_req_0 : boolean;
  signal phi_stmt_2448_req_1 : boolean;
  signal phi_stmt_2448_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeD_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeD_CP_5725_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeD_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_5725_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeD_CP_5725_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_5725_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeD_CP_5725: Block -- control-path 
    signal convTransposeD_CP_5725_elements: BooleanArray(91 downto 0);
    -- 
  begin -- 
    convTransposeD_CP_5725_elements(0) <= convTransposeD_CP_5725_start;
    convTransposeD_CP_5725_symbol <= convTransposeD_CP_5725_elements(67);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2299_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2299_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2299_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2297/$entry
      -- CP-element group 0: 	 branch_block_stmt_2297/branch_block_stmt_2297__entry__
      -- CP-element group 0: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333__entry__
      -- 
    rr_5773_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5773_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(0), ack => RPIPE_Block1_start_2299_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2299_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2299_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2299_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2299_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2299_update_start_
      -- CP-element group 1: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2299_sample_completed_
      -- 
    ra_5774_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2299_inst_ack_0, ack => convTransposeD_CP_5725_elements(1)); -- 
    cr_5778_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5778_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(1), ack => RPIPE_Block1_start_2299_inst_req_1); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2302_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2299_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2299_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2299_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2302_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2302_Sample/$entry
      -- 
    ca_5779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2299_inst_ack_1, ack => convTransposeD_CP_5725_elements(2)); -- 
    rr_5787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(2), ack => RPIPE_Block1_start_2302_inst_req_0); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2302_update_start_
      -- CP-element group 3: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2302_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2302_Update/cr
      -- CP-element group 3: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2302_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2302_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2302_Sample/$exit
      -- 
    ra_5788_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2302_inst_ack_0, ack => convTransposeD_CP_5725_elements(3)); -- 
    cr_5792_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5792_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(3), ack => RPIPE_Block1_start_2302_inst_req_1); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2302_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2305_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2302_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2305_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2302_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2305_Sample/rr
      -- 
    ca_5793_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2302_inst_ack_1, ack => convTransposeD_CP_5725_elements(4)); -- 
    rr_5801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(4), ack => RPIPE_Block1_start_2305_inst_req_0); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2305_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2305_update_start_
      -- CP-element group 5: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2305_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2305_Update/cr
      -- CP-element group 5: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2305_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2305_Update/$entry
      -- 
    ra_5802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2305_inst_ack_0, ack => convTransposeD_CP_5725_elements(5)); -- 
    cr_5806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(5), ack => RPIPE_Block1_start_2305_inst_req_1); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2305_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2308_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2305_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2308_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2305_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2308_sample_start_
      -- 
    ca_5807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2305_inst_ack_1, ack => convTransposeD_CP_5725_elements(6)); -- 
    rr_5815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(6), ack => RPIPE_Block1_start_2308_inst_req_0); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2308_Sample/ra
      -- CP-element group 7: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2308_Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2308_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2308_Update/cr
      -- CP-element group 7: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2308_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2308_update_start_
      -- 
    ra_5816_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2308_inst_ack_0, ack => convTransposeD_CP_5725_elements(7)); -- 
    cr_5820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(7), ack => RPIPE_Block1_start_2308_inst_req_1); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2308_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2311_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2311_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2308_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2308_Update/ca
      -- CP-element group 8: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2311_sample_start_
      -- 
    ca_5821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2308_inst_ack_1, ack => convTransposeD_CP_5725_elements(8)); -- 
    rr_5829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(8), ack => RPIPE_Block1_start_2311_inst_req_0); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2311_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2311_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2311_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2311_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2311_update_start_
      -- CP-element group 9: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2311_Update/cr
      -- 
    ra_5830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2311_inst_ack_0, ack => convTransposeD_CP_5725_elements(9)); -- 
    cr_5834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(9), ack => RPIPE_Block1_start_2311_inst_req_1); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2314_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2311_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2311_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2311_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2314_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2314_Sample/rr
      -- 
    ca_5835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2311_inst_ack_1, ack => convTransposeD_CP_5725_elements(10)); -- 
    rr_5843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(10), ack => RPIPE_Block1_start_2314_inst_req_0); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2314_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2314_update_start_
      -- CP-element group 11: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2314_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2314_Sample/ra
      -- CP-element group 11: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2314_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2314_Update/cr
      -- 
    ra_5844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2314_inst_ack_0, ack => convTransposeD_CP_5725_elements(11)); -- 
    cr_5848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(11), ack => RPIPE_Block1_start_2314_inst_req_1); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2314_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2314_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2314_Update/ca
      -- CP-element group 12: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2317_sample_start_
      -- CP-element group 12: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2317_Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2317_Sample/rr
      -- 
    ca_5849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2314_inst_ack_1, ack => convTransposeD_CP_5725_elements(12)); -- 
    rr_5857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(12), ack => RPIPE_Block1_start_2317_inst_req_0); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2317_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2317_update_start_
      -- CP-element group 13: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2317_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2317_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2317_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2317_Update/cr
      -- 
    ra_5858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2317_inst_ack_0, ack => convTransposeD_CP_5725_elements(13)); -- 
    cr_5862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(13), ack => RPIPE_Block1_start_2317_inst_req_1); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2317_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2317_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2317_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2320_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2320_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2320_Sample/rr
      -- 
    ca_5863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2317_inst_ack_1, ack => convTransposeD_CP_5725_elements(14)); -- 
    rr_5871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(14), ack => RPIPE_Block1_start_2320_inst_req_0); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2320_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2320_update_start_
      -- CP-element group 15: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2320_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2320_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2320_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2320_Update/cr
      -- 
    ra_5872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2320_inst_ack_0, ack => convTransposeD_CP_5725_elements(15)); -- 
    cr_5876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(15), ack => RPIPE_Block1_start_2320_inst_req_1); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2320_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2320_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2320_Update/ca
      -- CP-element group 16: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2323_sample_start_
      -- CP-element group 16: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2323_Sample/$entry
      -- CP-element group 16: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2323_Sample/rr
      -- 
    ca_5877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2320_inst_ack_1, ack => convTransposeD_CP_5725_elements(16)); -- 
    rr_5885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(16), ack => RPIPE_Block1_start_2323_inst_req_0); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2323_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2323_update_start_
      -- CP-element group 17: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2323_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2323_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2323_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2323_Update/cr
      -- 
    ra_5886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2323_inst_ack_0, ack => convTransposeD_CP_5725_elements(17)); -- 
    cr_5890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(17), ack => RPIPE_Block1_start_2323_inst_req_1); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2323_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2323_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2323_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2326_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2326_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2326_Sample/rr
      -- 
    ca_5891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2323_inst_ack_1, ack => convTransposeD_CP_5725_elements(18)); -- 
    rr_5899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(18), ack => RPIPE_Block1_start_2326_inst_req_0); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2326_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2326_update_start_
      -- CP-element group 19: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2326_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2326_Sample/ra
      -- CP-element group 19: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2326_Update/$entry
      -- CP-element group 19: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2326_Update/cr
      -- 
    ra_5900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2326_inst_ack_0, ack => convTransposeD_CP_5725_elements(19)); -- 
    cr_5904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(19), ack => RPIPE_Block1_start_2326_inst_req_1); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2326_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2326_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2326_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2329_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2329_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2329_Sample/rr
      -- 
    ca_5905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2326_inst_ack_1, ack => convTransposeD_CP_5725_elements(20)); -- 
    rr_5913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(20), ack => RPIPE_Block1_start_2329_inst_req_0); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2329_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2329_update_start_
      -- CP-element group 21: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2329_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2329_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2329_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2329_Update/cr
      -- 
    ra_5914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2329_inst_ack_0, ack => convTransposeD_CP_5725_elements(21)); -- 
    cr_5918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(21), ack => RPIPE_Block1_start_2329_inst_req_1); -- 
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (6) 
      -- CP-element group 22: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2329_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2329_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2329_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2332_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2332_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2332_Sample/rr
      -- 
    ca_5919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2329_inst_ack_1, ack => convTransposeD_CP_5725_elements(22)); -- 
    rr_5927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(22), ack => RPIPE_Block1_start_2332_inst_req_0); -- 
    -- CP-element group 23:  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (6) 
      -- CP-element group 23: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2332_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2332_update_start_
      -- CP-element group 23: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2332_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2332_Sample/ra
      -- CP-element group 23: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2332_Update/$entry
      -- CP-element group 23: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2332_Update/cr
      -- 
    ra_5928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2332_inst_ack_0, ack => convTransposeD_CP_5725_elements(23)); -- 
    cr_5932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(23), ack => RPIPE_Block1_start_2332_inst_req_1); -- 
    -- CP-element group 24:  fork  transition  place  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24: 	26 
    -- CP-element group 24: 	27 
    -- CP-element group 24: 	28 
    -- CP-element group 24: 	29 
    -- CP-element group 24: 	30 
    -- CP-element group 24:  members (25) 
      -- CP-element group 24: 	 branch_block_stmt_2297/assign_stmt_2340_to_assign_stmt_2380__entry__
      -- CP-element group 24: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/$exit
      -- CP-element group 24: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333__exit__
      -- CP-element group 24: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2332_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2332_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_2297/assign_stmt_2300_to_assign_stmt_2333/RPIPE_Block1_start_2332_Update/ca
      -- CP-element group 24: 	 branch_block_stmt_2297/assign_stmt_2340_to_assign_stmt_2380/$entry
      -- CP-element group 24: 	 branch_block_stmt_2297/assign_stmt_2340_to_assign_stmt_2380/type_cast_2349_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_2297/assign_stmt_2340_to_assign_stmt_2380/type_cast_2349_update_start_
      -- CP-element group 24: 	 branch_block_stmt_2297/assign_stmt_2340_to_assign_stmt_2380/type_cast_2349_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_2297/assign_stmt_2340_to_assign_stmt_2380/type_cast_2349_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_2297/assign_stmt_2340_to_assign_stmt_2380/type_cast_2349_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_2297/assign_stmt_2340_to_assign_stmt_2380/type_cast_2349_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_2297/assign_stmt_2340_to_assign_stmt_2380/type_cast_2353_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_2297/assign_stmt_2340_to_assign_stmt_2380/type_cast_2353_update_start_
      -- CP-element group 24: 	 branch_block_stmt_2297/assign_stmt_2340_to_assign_stmt_2380/type_cast_2353_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_2297/assign_stmt_2340_to_assign_stmt_2380/type_cast_2353_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_2297/assign_stmt_2340_to_assign_stmt_2380/type_cast_2353_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_2297/assign_stmt_2340_to_assign_stmt_2380/type_cast_2353_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_2297/assign_stmt_2340_to_assign_stmt_2380/type_cast_2357_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_2297/assign_stmt_2340_to_assign_stmt_2380/type_cast_2357_update_start_
      -- CP-element group 24: 	 branch_block_stmt_2297/assign_stmt_2340_to_assign_stmt_2380/type_cast_2357_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_2297/assign_stmt_2340_to_assign_stmt_2380/type_cast_2357_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_2297/assign_stmt_2340_to_assign_stmt_2380/type_cast_2357_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_2297/assign_stmt_2340_to_assign_stmt_2380/type_cast_2357_Update/cr
      -- 
    ca_5933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2332_inst_ack_1, ack => convTransposeD_CP_5725_elements(24)); -- 
    rr_5944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(24), ack => type_cast_2349_inst_req_0); -- 
    cr_5949_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5949_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(24), ack => type_cast_2349_inst_req_1); -- 
    rr_5958_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5958_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(24), ack => type_cast_2353_inst_req_0); -- 
    cr_5963_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5963_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(24), ack => type_cast_2353_inst_req_1); -- 
    rr_5972_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5972_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(24), ack => type_cast_2357_inst_req_0); -- 
    cr_5977_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5977_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(24), ack => type_cast_2357_inst_req_1); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_2297/assign_stmt_2340_to_assign_stmt_2380/type_cast_2349_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_2297/assign_stmt_2340_to_assign_stmt_2380/type_cast_2349_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_2297/assign_stmt_2340_to_assign_stmt_2380/type_cast_2349_Sample/ra
      -- 
    ra_5945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2349_inst_ack_0, ack => convTransposeD_CP_5725_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	31 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_2297/assign_stmt_2340_to_assign_stmt_2380/type_cast_2349_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_2297/assign_stmt_2340_to_assign_stmt_2380/type_cast_2349_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_2297/assign_stmt_2340_to_assign_stmt_2380/type_cast_2349_Update/ca
      -- 
    ca_5950_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2349_inst_ack_1, ack => convTransposeD_CP_5725_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	24 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_2297/assign_stmt_2340_to_assign_stmt_2380/type_cast_2353_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_2297/assign_stmt_2340_to_assign_stmt_2380/type_cast_2353_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_2297/assign_stmt_2340_to_assign_stmt_2380/type_cast_2353_Sample/ra
      -- 
    ra_5959_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2353_inst_ack_0, ack => convTransposeD_CP_5725_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	24 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	31 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_2297/assign_stmt_2340_to_assign_stmt_2380/type_cast_2353_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_2297/assign_stmt_2340_to_assign_stmt_2380/type_cast_2353_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_2297/assign_stmt_2340_to_assign_stmt_2380/type_cast_2353_Update/ca
      -- 
    ca_5964_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2353_inst_ack_1, ack => convTransposeD_CP_5725_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	24 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_2297/assign_stmt_2340_to_assign_stmt_2380/type_cast_2357_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_2297/assign_stmt_2340_to_assign_stmt_2380/type_cast_2357_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_2297/assign_stmt_2340_to_assign_stmt_2380/type_cast_2357_Sample/ra
      -- 
    ra_5973_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2357_inst_ack_0, ack => convTransposeD_CP_5725_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	24 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_2297/assign_stmt_2340_to_assign_stmt_2380/type_cast_2357_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_2297/assign_stmt_2340_to_assign_stmt_2380/type_cast_2357_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_2297/assign_stmt_2340_to_assign_stmt_2380/type_cast_2357_Update/ca
      -- 
    ca_5978_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2357_inst_ack_1, ack => convTransposeD_CP_5725_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  place  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	26 
    -- CP-element group 31: 	28 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	68 
    -- CP-element group 31: 	69 
    -- CP-element group 31: 	71 
    -- CP-element group 31: 	72 
    -- CP-element group 31:  members (20) 
      -- CP-element group 31: 	 branch_block_stmt_2297/entry_whilex_xbodyx_xouter
      -- CP-element group 31: 	 branch_block_stmt_2297/assign_stmt_2340_to_assign_stmt_2380__exit__
      -- CP-element group 31: 	 branch_block_stmt_2297/assign_stmt_2340_to_assign_stmt_2380/$exit
      -- CP-element group 31: 	 branch_block_stmt_2297/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 31: 	 branch_block_stmt_2297/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2383/$entry
      -- CP-element group 31: 	 branch_block_stmt_2297/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2383/phi_stmt_2383_sources/$entry
      -- CP-element group 31: 	 branch_block_stmt_2297/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2383/phi_stmt_2383_sources/type_cast_2386/$entry
      -- CP-element group 31: 	 branch_block_stmt_2297/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2383/phi_stmt_2383_sources/type_cast_2386/SplitProtocol/$entry
      -- CP-element group 31: 	 branch_block_stmt_2297/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2383/phi_stmt_2383_sources/type_cast_2386/SplitProtocol/Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2297/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2383/phi_stmt_2383_sources/type_cast_2386/SplitProtocol/Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_2297/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2383/phi_stmt_2383_sources/type_cast_2386/SplitProtocol/Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_2297/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2383/phi_stmt_2383_sources/type_cast_2386/SplitProtocol/Update/cr
      -- CP-element group 31: 	 branch_block_stmt_2297/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/$entry
      -- CP-element group 31: 	 branch_block_stmt_2297/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/$entry
      -- CP-element group 31: 	 branch_block_stmt_2297/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2394/$entry
      -- CP-element group 31: 	 branch_block_stmt_2297/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2394/SplitProtocol/$entry
      -- CP-element group 31: 	 branch_block_stmt_2297/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2394/SplitProtocol/Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2297/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2394/SplitProtocol/Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_2297/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2394/SplitProtocol/Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_2297/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2394/SplitProtocol/Update/cr
      -- 
    rr_6368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(31), ack => type_cast_2386_inst_req_0); -- 
    cr_6373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(31), ack => type_cast_2386_inst_req_1); -- 
    rr_6391_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6391_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(31), ack => type_cast_2394_inst_req_0); -- 
    cr_6396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(31), ack => type_cast_2394_inst_req_1); -- 
    convTransposeD_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_5725_elements(26) & convTransposeD_CP_5725_elements(28) & convTransposeD_CP_5725_elements(30);
      gj_convTransposeD_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_5725_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	91 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2475_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2475_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2475_Sample/ra
      -- 
    ra_5993_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2475_inst_ack_0, ack => convTransposeD_CP_5725_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	91 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2475_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2475_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2475_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2489_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2489_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2489_Sample/rr
      -- 
    ca_5998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2475_inst_ack_1, ack => convTransposeD_CP_5725_elements(33)); -- 
    rr_6006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(33), ack => type_cast_2489_inst_req_0); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2489_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2489_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2489_Sample/ra
      -- 
    ra_6007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2489_inst_ack_0, ack => convTransposeD_CP_5725_elements(34)); -- 
    -- CP-element group 35:  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	91 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (16) 
      -- CP-element group 35: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2489_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2489_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2489_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2495_index_resized_1
      -- CP-element group 35: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2495_index_scaled_1
      -- CP-element group 35: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2495_index_computed_1
      -- CP-element group 35: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2495_index_resize_1/$entry
      -- CP-element group 35: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2495_index_resize_1/$exit
      -- CP-element group 35: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2495_index_resize_1/index_resize_req
      -- CP-element group 35: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2495_index_resize_1/index_resize_ack
      -- CP-element group 35: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2495_index_scale_1/$entry
      -- CP-element group 35: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2495_index_scale_1/$exit
      -- CP-element group 35: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2495_index_scale_1/scale_rename_req
      -- CP-element group 35: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2495_index_scale_1/scale_rename_ack
      -- CP-element group 35: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2495_final_index_sum_regn_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2495_final_index_sum_regn_Sample/req
      -- 
    ca_6012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2489_inst_ack_1, ack => convTransposeD_CP_5725_elements(35)); -- 
    req_6037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(35), ack => array_obj_ref_2495_index_offset_req_0); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	55 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2495_final_index_sum_regn_sample_complete
      -- CP-element group 36: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2495_final_index_sum_regn_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2495_final_index_sum_regn_Sample/ack
      -- 
    ack_6038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2495_index_offset_ack_0, ack => convTransposeD_CP_5725_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	91 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (11) 
      -- CP-element group 37: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/addr_of_2496_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2495_root_address_calculated
      -- CP-element group 37: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2495_offset_calculated
      -- CP-element group 37: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2495_final_index_sum_regn_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2495_final_index_sum_regn_Update/ack
      -- CP-element group 37: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2495_base_plus_offset/$entry
      -- CP-element group 37: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2495_base_plus_offset/$exit
      -- CP-element group 37: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2495_base_plus_offset/sum_rename_req
      -- CP-element group 37: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2495_base_plus_offset/sum_rename_ack
      -- CP-element group 37: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/addr_of_2496_request/$entry
      -- CP-element group 37: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/addr_of_2496_request/req
      -- 
    ack_6043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2495_index_offset_ack_1, ack => convTransposeD_CP_5725_elements(37)); -- 
    req_6052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(37), ack => addr_of_2496_final_reg_req_0); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/addr_of_2496_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/addr_of_2496_request/$exit
      -- CP-element group 38: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/addr_of_2496_request/ack
      -- 
    ack_6053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2496_final_reg_ack_0, ack => convTransposeD_CP_5725_elements(38)); -- 
    -- CP-element group 39:  join  fork  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	91 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (24) 
      -- CP-element group 39: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/addr_of_2496_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/addr_of_2496_complete/$exit
      -- CP-element group 39: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/addr_of_2496_complete/ack
      -- CP-element group 39: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2500_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2500_base_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2500_word_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2500_root_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2500_base_address_resized
      -- CP-element group 39: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2500_base_addr_resize/$entry
      -- CP-element group 39: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2500_base_addr_resize/$exit
      -- CP-element group 39: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2500_base_addr_resize/base_resize_req
      -- CP-element group 39: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2500_base_addr_resize/base_resize_ack
      -- CP-element group 39: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2500_base_plus_offset/$entry
      -- CP-element group 39: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2500_base_plus_offset/$exit
      -- CP-element group 39: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2500_base_plus_offset/sum_rename_req
      -- CP-element group 39: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2500_base_plus_offset/sum_rename_ack
      -- CP-element group 39: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2500_word_addrgen/$entry
      -- CP-element group 39: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2500_word_addrgen/$exit
      -- CP-element group 39: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2500_word_addrgen/root_register_req
      -- CP-element group 39: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2500_word_addrgen/root_register_ack
      -- CP-element group 39: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2500_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2500_Sample/word_access_start/$entry
      -- CP-element group 39: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2500_Sample/word_access_start/word_0/$entry
      -- CP-element group 39: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2500_Sample/word_access_start/word_0/rr
      -- 
    ack_6058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2496_final_reg_ack_1, ack => convTransposeD_CP_5725_elements(39)); -- 
    rr_6091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(39), ack => ptr_deref_2500_load_0_req_0); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (5) 
      -- CP-element group 40: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2500_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2500_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2500_Sample/word_access_start/$exit
      -- CP-element group 40: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2500_Sample/word_access_start/word_0/$exit
      -- CP-element group 40: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2500_Sample/word_access_start/word_0/ra
      -- 
    ra_6092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2500_load_0_ack_0, ack => convTransposeD_CP_5725_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	91 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	50 
    -- CP-element group 41:  members (9) 
      -- CP-element group 41: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2500_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2500_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2500_Update/word_access_complete/$exit
      -- CP-element group 41: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2500_Update/word_access_complete/word_0/$exit
      -- CP-element group 41: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2500_Update/word_access_complete/word_0/ca
      -- CP-element group 41: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2500_Update/ptr_deref_2500_Merge/$entry
      -- CP-element group 41: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2500_Update/ptr_deref_2500_Merge/$exit
      -- CP-element group 41: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2500_Update/ptr_deref_2500_Merge/merge_req
      -- CP-element group 41: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2500_Update/ptr_deref_2500_Merge/merge_ack
      -- 
    ca_6103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2500_load_0_ack_1, ack => convTransposeD_CP_5725_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	91 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2505_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2505_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2505_Sample/ra
      -- 
    ra_6117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2505_inst_ack_0, ack => convTransposeD_CP_5725_elements(42)); -- 
    -- CP-element group 43:  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	91 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (6) 
      -- CP-element group 43: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2505_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2505_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2505_Update/ca
      -- CP-element group 43: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2519_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2519_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2519_Sample/rr
      -- 
    ca_6122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2505_inst_ack_1, ack => convTransposeD_CP_5725_elements(43)); -- 
    rr_6130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(43), ack => type_cast_2519_inst_req_0); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2519_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2519_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2519_Sample/ra
      -- 
    ra_6131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2519_inst_ack_0, ack => convTransposeD_CP_5725_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	91 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (16) 
      -- CP-element group 45: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2519_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2519_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2519_Update/ca
      -- CP-element group 45: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2525_index_resized_1
      -- CP-element group 45: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2525_index_scaled_1
      -- CP-element group 45: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2525_index_computed_1
      -- CP-element group 45: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2525_index_resize_1/$entry
      -- CP-element group 45: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2525_index_resize_1/$exit
      -- CP-element group 45: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2525_index_resize_1/index_resize_req
      -- CP-element group 45: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2525_index_resize_1/index_resize_ack
      -- CP-element group 45: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2525_index_scale_1/$entry
      -- CP-element group 45: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2525_index_scale_1/$exit
      -- CP-element group 45: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2525_index_scale_1/scale_rename_req
      -- CP-element group 45: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2525_index_scale_1/scale_rename_ack
      -- CP-element group 45: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2525_final_index_sum_regn_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2525_final_index_sum_regn_Sample/req
      -- 
    ca_6136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2519_inst_ack_1, ack => convTransposeD_CP_5725_elements(45)); -- 
    req_6161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(45), ack => array_obj_ref_2525_index_offset_req_0); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	55 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2525_final_index_sum_regn_sample_complete
      -- CP-element group 46: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2525_final_index_sum_regn_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2525_final_index_sum_regn_Sample/ack
      -- 
    ack_6162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2525_index_offset_ack_0, ack => convTransposeD_CP_5725_elements(46)); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	91 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (11) 
      -- CP-element group 47: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/addr_of_2526_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2525_root_address_calculated
      -- CP-element group 47: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2525_offset_calculated
      -- CP-element group 47: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2525_final_index_sum_regn_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2525_final_index_sum_regn_Update/ack
      -- CP-element group 47: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2525_base_plus_offset/$entry
      -- CP-element group 47: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2525_base_plus_offset/$exit
      -- CP-element group 47: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2525_base_plus_offset/sum_rename_req
      -- CP-element group 47: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2525_base_plus_offset/sum_rename_ack
      -- CP-element group 47: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/addr_of_2526_request/$entry
      -- CP-element group 47: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/addr_of_2526_request/req
      -- 
    ack_6167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2525_index_offset_ack_1, ack => convTransposeD_CP_5725_elements(47)); -- 
    req_6176_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6176_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(47), ack => addr_of_2526_final_reg_req_0); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/addr_of_2526_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/addr_of_2526_request/$exit
      -- CP-element group 48: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/addr_of_2526_request/ack
      -- 
    ack_6177_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2526_final_reg_ack_0, ack => convTransposeD_CP_5725_elements(48)); -- 
    -- CP-element group 49:  fork  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	91 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (19) 
      -- CP-element group 49: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/addr_of_2526_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/addr_of_2526_complete/$exit
      -- CP-element group 49: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/addr_of_2526_complete/ack
      -- CP-element group 49: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2529_base_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2529_word_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2529_root_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2529_base_address_resized
      -- CP-element group 49: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2529_base_addr_resize/$entry
      -- CP-element group 49: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2529_base_addr_resize/$exit
      -- CP-element group 49: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2529_base_addr_resize/base_resize_req
      -- CP-element group 49: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2529_base_addr_resize/base_resize_ack
      -- CP-element group 49: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2529_base_plus_offset/$entry
      -- CP-element group 49: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2529_base_plus_offset/$exit
      -- CP-element group 49: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2529_base_plus_offset/sum_rename_req
      -- CP-element group 49: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2529_base_plus_offset/sum_rename_ack
      -- CP-element group 49: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2529_word_addrgen/$entry
      -- CP-element group 49: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2529_word_addrgen/$exit
      -- CP-element group 49: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2529_word_addrgen/root_register_req
      -- CP-element group 49: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2529_word_addrgen/root_register_ack
      -- 
    ack_6182_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2526_final_reg_ack_1, ack => convTransposeD_CP_5725_elements(49)); -- 
    -- CP-element group 50:  join  transition  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	41 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2529_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2529_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2529_Sample/ptr_deref_2529_Split/$entry
      -- CP-element group 50: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2529_Sample/ptr_deref_2529_Split/$exit
      -- CP-element group 50: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2529_Sample/ptr_deref_2529_Split/split_req
      -- CP-element group 50: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2529_Sample/ptr_deref_2529_Split/split_ack
      -- CP-element group 50: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2529_Sample/word_access_start/$entry
      -- CP-element group 50: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2529_Sample/word_access_start/word_0/$entry
      -- CP-element group 50: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2529_Sample/word_access_start/word_0/rr
      -- 
    rr_6220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(50), ack => ptr_deref_2529_store_0_req_0); -- 
    convTransposeD_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_5725_elements(41) & convTransposeD_CP_5725_elements(49);
      gj_convTransposeD_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_5725_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (5) 
      -- CP-element group 51: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2529_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2529_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2529_Sample/word_access_start/$exit
      -- CP-element group 51: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2529_Sample/word_access_start/word_0/$exit
      -- CP-element group 51: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2529_Sample/word_access_start/word_0/ra
      -- 
    ra_6221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2529_store_0_ack_0, ack => convTransposeD_CP_5725_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	91 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	55 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2529_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2529_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2529_Update/word_access_complete/$exit
      -- CP-element group 52: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2529_Update/word_access_complete/word_0/$exit
      -- CP-element group 52: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2529_Update/word_access_complete/word_0/ca
      -- 
    ca_6232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2529_store_0_ack_1, ack => convTransposeD_CP_5725_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	91 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2535_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2535_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2535_Sample/ra
      -- 
    ra_6241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2535_inst_ack_0, ack => convTransposeD_CP_5725_elements(53)); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	91 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2535_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2535_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2535_Update/ca
      -- 
    ca_6246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2535_inst_ack_1, ack => convTransposeD_CP_5725_elements(54)); -- 
    -- CP-element group 55:  branch  join  transition  place  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	36 
    -- CP-element group 55: 	46 
    -- CP-element group 55: 	52 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (10) 
      -- CP-element group 55: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549__exit__
      -- CP-element group 55: 	 branch_block_stmt_2297/if_stmt_2550__entry__
      -- CP-element group 55: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/$exit
      -- CP-element group 55: 	 branch_block_stmt_2297/if_stmt_2550_dead_link/$entry
      -- CP-element group 55: 	 branch_block_stmt_2297/if_stmt_2550_eval_test/$entry
      -- CP-element group 55: 	 branch_block_stmt_2297/if_stmt_2550_eval_test/$exit
      -- CP-element group 55: 	 branch_block_stmt_2297/if_stmt_2550_eval_test/branch_req
      -- CP-element group 55: 	 branch_block_stmt_2297/R_cmp_2551_place
      -- CP-element group 55: 	 branch_block_stmt_2297/if_stmt_2550_if_link/$entry
      -- CP-element group 55: 	 branch_block_stmt_2297/if_stmt_2550_else_link/$entry
      -- 
    branch_req_6254_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6254_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(55), ack => if_stmt_2550_branch_req_0); -- 
    convTransposeD_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_5725_elements(36) & convTransposeD_CP_5725_elements(46) & convTransposeD_CP_5725_elements(52) & convTransposeD_CP_5725_elements(54);
      gj_convTransposeD_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_5725_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	86 
    -- CP-element group 56: 	87 
    -- CP-element group 56:  members (24) 
      -- CP-element group 56: 	 branch_block_stmt_2297/assign_stmt_2562__entry__
      -- CP-element group 56: 	 branch_block_stmt_2297/ifx_xthen_whilex_xbody
      -- CP-element group 56: 	 branch_block_stmt_2297/assign_stmt_2562__exit__
      -- CP-element group 56: 	 branch_block_stmt_2297/merge_stmt_2556__exit__
      -- CP-element group 56: 	 branch_block_stmt_2297/if_stmt_2550_if_link/$exit
      -- CP-element group 56: 	 branch_block_stmt_2297/if_stmt_2550_if_link/if_choice_transition
      -- CP-element group 56: 	 branch_block_stmt_2297/whilex_xbody_ifx_xthen
      -- CP-element group 56: 	 branch_block_stmt_2297/assign_stmt_2562/$entry
      -- CP-element group 56: 	 branch_block_stmt_2297/assign_stmt_2562/$exit
      -- CP-element group 56: 	 branch_block_stmt_2297/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 56: 	 branch_block_stmt_2297/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2448/$entry
      -- CP-element group 56: 	 branch_block_stmt_2297/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/$entry
      -- CP-element group 56: 	 branch_block_stmt_2297/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/type_cast_2451/$entry
      -- CP-element group 56: 	 branch_block_stmt_2297/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/type_cast_2451/SplitProtocol/$entry
      -- CP-element group 56: 	 branch_block_stmt_2297/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/type_cast_2451/SplitProtocol/Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_2297/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/type_cast_2451/SplitProtocol/Sample/rr
      -- CP-element group 56: 	 branch_block_stmt_2297/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/type_cast_2451/SplitProtocol/Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_2297/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/type_cast_2451/SplitProtocol/Update/cr
      -- CP-element group 56: 	 branch_block_stmt_2297/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 56: 	 branch_block_stmt_2297/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 56: 	 branch_block_stmt_2297/merge_stmt_2556_PhiReqMerge
      -- CP-element group 56: 	 branch_block_stmt_2297/merge_stmt_2556_PhiAck/$entry
      -- CP-element group 56: 	 branch_block_stmt_2297/merge_stmt_2556_PhiAck/$exit
      -- CP-element group 56: 	 branch_block_stmt_2297/merge_stmt_2556_PhiAck/dummy
      -- 
    if_choice_transition_6259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2550_branch_ack_1, ack => convTransposeD_CP_5725_elements(56)); -- 
    rr_6472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(56), ack => type_cast_2451_inst_req_0); -- 
    cr_6477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(56), ack => type_cast_2451_inst_req_1); -- 
    -- CP-element group 57:  fork  transition  place  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57: 	59 
    -- CP-element group 57: 	61 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (24) 
      -- CP-element group 57: 	 branch_block_stmt_2297/merge_stmt_2564__exit__
      -- CP-element group 57: 	 branch_block_stmt_2297/assign_stmt_2570_to_assign_stmt_2605__entry__
      -- CP-element group 57: 	 branch_block_stmt_2297/if_stmt_2550_else_link/$exit
      -- CP-element group 57: 	 branch_block_stmt_2297/if_stmt_2550_else_link/else_choice_transition
      -- CP-element group 57: 	 branch_block_stmt_2297/whilex_xbody_ifx_xelse
      -- CP-element group 57: 	 branch_block_stmt_2297/assign_stmt_2570_to_assign_stmt_2605/$entry
      -- CP-element group 57: 	 branch_block_stmt_2297/assign_stmt_2570_to_assign_stmt_2605/type_cast_2574_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_2297/assign_stmt_2570_to_assign_stmt_2605/type_cast_2574_update_start_
      -- CP-element group 57: 	 branch_block_stmt_2297/merge_stmt_2564_PhiReqMerge
      -- CP-element group 57: 	 branch_block_stmt_2297/assign_stmt_2570_to_assign_stmt_2605/type_cast_2574_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_2297/assign_stmt_2570_to_assign_stmt_2605/type_cast_2574_Sample/rr
      -- CP-element group 57: 	 branch_block_stmt_2297/merge_stmt_2564_PhiAck/dummy
      -- CP-element group 57: 	 branch_block_stmt_2297/assign_stmt_2570_to_assign_stmt_2605/type_cast_2574_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_2297/assign_stmt_2570_to_assign_stmt_2605/type_cast_2574_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_2297/assign_stmt_2570_to_assign_stmt_2605/type_cast_2589_update_start_
      -- CP-element group 57: 	 branch_block_stmt_2297/merge_stmt_2564_PhiAck/$exit
      -- CP-element group 57: 	 branch_block_stmt_2297/assign_stmt_2570_to_assign_stmt_2605/type_cast_2589_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_2297/assign_stmt_2570_to_assign_stmt_2605/type_cast_2589_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_2297/assign_stmt_2570_to_assign_stmt_2605/type_cast_2599_update_start_
      -- CP-element group 57: 	 branch_block_stmt_2297/merge_stmt_2564_PhiAck/$entry
      -- CP-element group 57: 	 branch_block_stmt_2297/assign_stmt_2570_to_assign_stmt_2605/type_cast_2599_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_2297/assign_stmt_2570_to_assign_stmt_2605/type_cast_2599_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_2297/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 57: 	 branch_block_stmt_2297/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- 
    else_choice_transition_6263_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2550_branch_ack_0, ack => convTransposeD_CP_5725_elements(57)); -- 
    rr_6279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(57), ack => type_cast_2574_inst_req_0); -- 
    cr_6284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(57), ack => type_cast_2574_inst_req_1); -- 
    cr_6298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(57), ack => type_cast_2589_inst_req_1); -- 
    cr_6312_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6312_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(57), ack => type_cast_2599_inst_req_1); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_2297/assign_stmt_2570_to_assign_stmt_2605/type_cast_2574_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_2297/assign_stmt_2570_to_assign_stmt_2605/type_cast_2574_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_2297/assign_stmt_2570_to_assign_stmt_2605/type_cast_2574_Sample/ra
      -- 
    ra_6280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2574_inst_ack_0, ack => convTransposeD_CP_5725_elements(58)); -- 
    -- CP-element group 59:  transition  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (6) 
      -- CP-element group 59: 	 branch_block_stmt_2297/assign_stmt_2570_to_assign_stmt_2605/type_cast_2574_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_2297/assign_stmt_2570_to_assign_stmt_2605/type_cast_2574_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_2297/assign_stmt_2570_to_assign_stmt_2605/type_cast_2574_Update/ca
      -- CP-element group 59: 	 branch_block_stmt_2297/assign_stmt_2570_to_assign_stmt_2605/type_cast_2589_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_2297/assign_stmt_2570_to_assign_stmt_2605/type_cast_2589_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_2297/assign_stmt_2570_to_assign_stmt_2605/type_cast_2589_Sample/rr
      -- 
    ca_6285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2574_inst_ack_1, ack => convTransposeD_CP_5725_elements(59)); -- 
    rr_6293_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6293_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(59), ack => type_cast_2589_inst_req_0); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_2297/assign_stmt_2570_to_assign_stmt_2605/type_cast_2589_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_2297/assign_stmt_2570_to_assign_stmt_2605/type_cast_2589_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_2297/assign_stmt_2570_to_assign_stmt_2605/type_cast_2589_Sample/ra
      -- 
    ra_6294_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2589_inst_ack_0, ack => convTransposeD_CP_5725_elements(60)); -- 
    -- CP-element group 61:  transition  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	57 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_2297/assign_stmt_2570_to_assign_stmt_2605/type_cast_2589_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_2297/assign_stmt_2570_to_assign_stmt_2605/type_cast_2589_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_2297/assign_stmt_2570_to_assign_stmt_2605/type_cast_2589_Update/ca
      -- CP-element group 61: 	 branch_block_stmt_2297/assign_stmt_2570_to_assign_stmt_2605/type_cast_2599_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_2297/assign_stmt_2570_to_assign_stmt_2605/type_cast_2599_Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_2297/assign_stmt_2570_to_assign_stmt_2605/type_cast_2599_Sample/rr
      -- 
    ca_6299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2589_inst_ack_1, ack => convTransposeD_CP_5725_elements(61)); -- 
    rr_6307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(61), ack => type_cast_2599_inst_req_0); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_2297/assign_stmt_2570_to_assign_stmt_2605/type_cast_2599_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_2297/assign_stmt_2570_to_assign_stmt_2605/type_cast_2599_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_2297/assign_stmt_2570_to_assign_stmt_2605/type_cast_2599_Sample/ra
      -- 
    ra_6308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2599_inst_ack_0, ack => convTransposeD_CP_5725_elements(62)); -- 
    -- CP-element group 63:  branch  transition  place  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (13) 
      -- CP-element group 63: 	 branch_block_stmt_2297/assign_stmt_2570_to_assign_stmt_2605__exit__
      -- CP-element group 63: 	 branch_block_stmt_2297/if_stmt_2606__entry__
      -- CP-element group 63: 	 branch_block_stmt_2297/assign_stmt_2570_to_assign_stmt_2605/$exit
      -- CP-element group 63: 	 branch_block_stmt_2297/assign_stmt_2570_to_assign_stmt_2605/type_cast_2599_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_2297/assign_stmt_2570_to_assign_stmt_2605/type_cast_2599_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_2297/assign_stmt_2570_to_assign_stmt_2605/type_cast_2599_Update/ca
      -- CP-element group 63: 	 branch_block_stmt_2297/if_stmt_2606_dead_link/$entry
      -- CP-element group 63: 	 branch_block_stmt_2297/if_stmt_2606_eval_test/$entry
      -- CP-element group 63: 	 branch_block_stmt_2297/if_stmt_2606_eval_test/$exit
      -- CP-element group 63: 	 branch_block_stmt_2297/if_stmt_2606_eval_test/branch_req
      -- CP-element group 63: 	 branch_block_stmt_2297/R_cmp137_2607_place
      -- CP-element group 63: 	 branch_block_stmt_2297/if_stmt_2606_if_link/$entry
      -- CP-element group 63: 	 branch_block_stmt_2297/if_stmt_2606_else_link/$entry
      -- 
    ca_6313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2599_inst_ack_1, ack => convTransposeD_CP_5725_elements(63)); -- 
    branch_req_6321_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6321_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(63), ack => if_stmt_2606_branch_req_0); -- 
    -- CP-element group 64:  merge  transition  place  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (15) 
      -- CP-element group 64: 	 branch_block_stmt_2297/assign_stmt_2617__entry__
      -- CP-element group 64: 	 branch_block_stmt_2297/merge_stmt_2612__exit__
      -- CP-element group 64: 	 branch_block_stmt_2297/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 64: 	 branch_block_stmt_2297/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 64: 	 branch_block_stmt_2297/merge_stmt_2612_PhiAck/$entry
      -- CP-element group 64: 	 branch_block_stmt_2297/merge_stmt_2612_PhiAck/$exit
      -- CP-element group 64: 	 branch_block_stmt_2297/merge_stmt_2612_PhiAck/dummy
      -- CP-element group 64: 	 branch_block_stmt_2297/merge_stmt_2612_PhiReqMerge
      -- CP-element group 64: 	 branch_block_stmt_2297/if_stmt_2606_if_link/$exit
      -- CP-element group 64: 	 branch_block_stmt_2297/if_stmt_2606_if_link/if_choice_transition
      -- CP-element group 64: 	 branch_block_stmt_2297/ifx_xelse_whilex_xend
      -- CP-element group 64: 	 branch_block_stmt_2297/assign_stmt_2617/$entry
      -- CP-element group 64: 	 branch_block_stmt_2297/assign_stmt_2617/WPIPE_Block3_done_2614_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_2297/assign_stmt_2617/WPIPE_Block3_done_2614_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_2297/assign_stmt_2617/WPIPE_Block3_done_2614_Sample/req
      -- 
    if_choice_transition_6326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2606_branch_ack_1, ack => convTransposeD_CP_5725_elements(64)); -- 
    req_6343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(64), ack => WPIPE_Block3_done_2614_inst_req_0); -- 
    -- CP-element group 65:  fork  transition  place  input  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	75 
    -- CP-element group 65: 	76 
    -- CP-element group 65: 	78 
    -- CP-element group 65: 	79 
    -- CP-element group 65:  members (20) 
      -- CP-element group 65: 	 branch_block_stmt_2297/if_stmt_2606_else_link/$exit
      -- CP-element group 65: 	 branch_block_stmt_2297/if_stmt_2606_else_link/else_choice_transition
      -- CP-element group 65: 	 branch_block_stmt_2297/ifx_xelse_whilex_xbodyx_xouter
      -- CP-element group 65: 	 branch_block_stmt_2297/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 65: 	 branch_block_stmt_2297/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2383/$entry
      -- CP-element group 65: 	 branch_block_stmt_2297/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2383/phi_stmt_2383_sources/$entry
      -- CP-element group 65: 	 branch_block_stmt_2297/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2383/phi_stmt_2383_sources/type_cast_2388/$entry
      -- CP-element group 65: 	 branch_block_stmt_2297/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2383/phi_stmt_2383_sources/type_cast_2388/SplitProtocol/$entry
      -- CP-element group 65: 	 branch_block_stmt_2297/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2383/phi_stmt_2383_sources/type_cast_2388/SplitProtocol/Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_2297/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2383/phi_stmt_2383_sources/type_cast_2388/SplitProtocol/Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_2297/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2383/phi_stmt_2383_sources/type_cast_2388/SplitProtocol/Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_2297/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2383/phi_stmt_2383_sources/type_cast_2388/SplitProtocol/Update/cr
      -- CP-element group 65: 	 branch_block_stmt_2297/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/$entry
      -- CP-element group 65: 	 branch_block_stmt_2297/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/$entry
      -- CP-element group 65: 	 branch_block_stmt_2297/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2392/$entry
      -- CP-element group 65: 	 branch_block_stmt_2297/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2392/SplitProtocol/$entry
      -- CP-element group 65: 	 branch_block_stmt_2297/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2392/SplitProtocol/Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_2297/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2392/SplitProtocol/Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_2297/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2392/SplitProtocol/Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_2297/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2392/SplitProtocol/Update/cr
      -- 
    else_choice_transition_6330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2606_branch_ack_0, ack => convTransposeD_CP_5725_elements(65)); -- 
    rr_6417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(65), ack => type_cast_2388_inst_req_0); -- 
    cr_6422_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6422_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(65), ack => type_cast_2388_inst_req_1); -- 
    rr_6440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(65), ack => type_cast_2392_inst_req_0); -- 
    cr_6445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(65), ack => type_cast_2392_inst_req_1); -- 
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_2297/assign_stmt_2617/WPIPE_Block3_done_2614_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_2297/assign_stmt_2617/WPIPE_Block3_done_2614_update_start_
      -- CP-element group 66: 	 branch_block_stmt_2297/assign_stmt_2617/WPIPE_Block3_done_2614_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_2297/assign_stmt_2617/WPIPE_Block3_done_2614_Sample/ack
      -- CP-element group 66: 	 branch_block_stmt_2297/assign_stmt_2617/WPIPE_Block3_done_2614_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_2297/assign_stmt_2617/WPIPE_Block3_done_2614_Update/req
      -- 
    ack_6344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_2614_inst_ack_0, ack => convTransposeD_CP_5725_elements(66)); -- 
    req_6348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(66), ack => WPIPE_Block3_done_2614_inst_req_1); -- 
    -- CP-element group 67:  transition  place  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (16) 
      -- CP-element group 67: 	 branch_block_stmt_2297/merge_stmt_2619__exit__
      -- CP-element group 67: 	 branch_block_stmt_2297/return__
      -- CP-element group 67: 	 branch_block_stmt_2297/assign_stmt_2617__exit__
      -- CP-element group 67: 	 branch_block_stmt_2297/merge_stmt_2619_PhiReqMerge
      -- CP-element group 67: 	 branch_block_stmt_2297/return___PhiReq/$entry
      -- CP-element group 67: 	 branch_block_stmt_2297/return___PhiReq/$exit
      -- CP-element group 67: 	 $exit
      -- CP-element group 67: 	 branch_block_stmt_2297/$exit
      -- CP-element group 67: 	 branch_block_stmt_2297/branch_block_stmt_2297__exit__
      -- CP-element group 67: 	 branch_block_stmt_2297/assign_stmt_2617/$exit
      -- CP-element group 67: 	 branch_block_stmt_2297/assign_stmt_2617/WPIPE_Block3_done_2614_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_2297/assign_stmt_2617/WPIPE_Block3_done_2614_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_2297/assign_stmt_2617/WPIPE_Block3_done_2614_Update/ack
      -- CP-element group 67: 	 branch_block_stmt_2297/merge_stmt_2619_PhiAck/dummy
      -- CP-element group 67: 	 branch_block_stmt_2297/merge_stmt_2619_PhiAck/$exit
      -- CP-element group 67: 	 branch_block_stmt_2297/merge_stmt_2619_PhiAck/$entry
      -- 
    ack_6349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_2614_inst_ack_1, ack => convTransposeD_CP_5725_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	31 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (2) 
      -- CP-element group 68: 	 branch_block_stmt_2297/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2383/phi_stmt_2383_sources/type_cast_2386/SplitProtocol/Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_2297/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2383/phi_stmt_2383_sources/type_cast_2386/SplitProtocol/Sample/ra
      -- 
    ra_6369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2386_inst_ack_0, ack => convTransposeD_CP_5725_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	31 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (2) 
      -- CP-element group 69: 	 branch_block_stmt_2297/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2383/phi_stmt_2383_sources/type_cast_2386/SplitProtocol/Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_2297/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2383/phi_stmt_2383_sources/type_cast_2386/SplitProtocol/Update/ca
      -- 
    ca_6374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2386_inst_ack_1, ack => convTransposeD_CP_5725_elements(69)); -- 
    -- CP-element group 70:  join  transition  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	74 
    -- CP-element group 70:  members (5) 
      -- CP-element group 70: 	 branch_block_stmt_2297/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2383/$exit
      -- CP-element group 70: 	 branch_block_stmt_2297/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2383/phi_stmt_2383_sources/$exit
      -- CP-element group 70: 	 branch_block_stmt_2297/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2383/phi_stmt_2383_sources/type_cast_2386/$exit
      -- CP-element group 70: 	 branch_block_stmt_2297/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2383/phi_stmt_2383_sources/type_cast_2386/SplitProtocol/$exit
      -- CP-element group 70: 	 branch_block_stmt_2297/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2383/phi_stmt_2383_req
      -- 
    phi_stmt_2383_req_6375_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2383_req_6375_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(70), ack => phi_stmt_2383_req_0); -- 
    convTransposeD_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_5725_elements(68) & convTransposeD_CP_5725_elements(69);
      gj_convTransposeD_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_5725_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	31 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (2) 
      -- CP-element group 71: 	 branch_block_stmt_2297/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2394/SplitProtocol/Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_2297/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2394/SplitProtocol/Sample/ra
      -- 
    ra_6392_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2394_inst_ack_0, ack => convTransposeD_CP_5725_elements(71)); -- 
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	31 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (2) 
      -- CP-element group 72: 	 branch_block_stmt_2297/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2394/SplitProtocol/Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_2297/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2394/SplitProtocol/Update/ca
      -- 
    ca_6397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2394_inst_ack_1, ack => convTransposeD_CP_5725_elements(72)); -- 
    -- CP-element group 73:  join  transition  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (5) 
      -- CP-element group 73: 	 branch_block_stmt_2297/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/$exit
      -- CP-element group 73: 	 branch_block_stmt_2297/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/$exit
      -- CP-element group 73: 	 branch_block_stmt_2297/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2394/$exit
      -- CP-element group 73: 	 branch_block_stmt_2297/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2394/SplitProtocol/$exit
      -- CP-element group 73: 	 branch_block_stmt_2297/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_req
      -- 
    phi_stmt_2389_req_6398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2389_req_6398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(73), ack => phi_stmt_2389_req_1); -- 
    convTransposeD_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_5725_elements(71) & convTransposeD_CP_5725_elements(72);
      gj_convTransposeD_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_5725_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  join  transition  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	70 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	82 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_2297/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_5725_elements(70) & convTransposeD_CP_5725_elements(73);
      gj_convTransposeD_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_5725_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	65 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_2297/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2383/phi_stmt_2383_sources/type_cast_2388/SplitProtocol/Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_2297/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2383/phi_stmt_2383_sources/type_cast_2388/SplitProtocol/Sample/ra
      -- 
    ra_6418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2388_inst_ack_0, ack => convTransposeD_CP_5725_elements(75)); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	65 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (2) 
      -- CP-element group 76: 	 branch_block_stmt_2297/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2383/phi_stmt_2383_sources/type_cast_2388/SplitProtocol/Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_2297/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2383/phi_stmt_2383_sources/type_cast_2388/SplitProtocol/Update/ca
      -- 
    ca_6423_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2388_inst_ack_1, ack => convTransposeD_CP_5725_elements(76)); -- 
    -- CP-element group 77:  join  transition  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	81 
    -- CP-element group 77:  members (5) 
      -- CP-element group 77: 	 branch_block_stmt_2297/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2383/$exit
      -- CP-element group 77: 	 branch_block_stmt_2297/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2383/phi_stmt_2383_sources/$exit
      -- CP-element group 77: 	 branch_block_stmt_2297/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2383/phi_stmt_2383_sources/type_cast_2388/$exit
      -- CP-element group 77: 	 branch_block_stmt_2297/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2383/phi_stmt_2383_sources/type_cast_2388/SplitProtocol/$exit
      -- CP-element group 77: 	 branch_block_stmt_2297/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2383/phi_stmt_2383_req
      -- 
    phi_stmt_2383_req_6424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2383_req_6424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(77), ack => phi_stmt_2383_req_1); -- 
    convTransposeD_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_5725_elements(75) & convTransposeD_CP_5725_elements(76);
      gj_convTransposeD_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_5725_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	65 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (2) 
      -- CP-element group 78: 	 branch_block_stmt_2297/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2392/SplitProtocol/Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_2297/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2392/SplitProtocol/Sample/ra
      -- 
    ra_6441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2392_inst_ack_0, ack => convTransposeD_CP_5725_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	65 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_2297/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2392/SplitProtocol/Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_2297/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2392/SplitProtocol/Update/ca
      -- 
    ca_6446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2392_inst_ack_1, ack => convTransposeD_CP_5725_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (5) 
      -- CP-element group 80: 	 branch_block_stmt_2297/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/$exit
      -- CP-element group 80: 	 branch_block_stmt_2297/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/$exit
      -- CP-element group 80: 	 branch_block_stmt_2297/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2392/$exit
      -- CP-element group 80: 	 branch_block_stmt_2297/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2392/SplitProtocol/$exit
      -- CP-element group 80: 	 branch_block_stmt_2297/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_req
      -- 
    phi_stmt_2389_req_6447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2389_req_6447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(80), ack => phi_stmt_2389_req_0); -- 
    convTransposeD_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_5725_elements(78) & convTransposeD_CP_5725_elements(79);
      gj_convTransposeD_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_5725_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  join  transition  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	77 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_2297/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_5725_elements(77) & convTransposeD_CP_5725_elements(80);
      gj_convTransposeD_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_5725_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  merge  fork  transition  place  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	74 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_2297/merge_stmt_2382_PhiReqMerge
      -- CP-element group 82: 	 branch_block_stmt_2297/merge_stmt_2382_PhiAck/$entry
      -- 
    convTransposeD_CP_5725_elements(82) <= OrReduce(convTransposeD_CP_5725_elements(74) & convTransposeD_CP_5725_elements(81));
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (1) 
      -- CP-element group 83: 	 branch_block_stmt_2297/merge_stmt_2382_PhiAck/phi_stmt_2383_ack
      -- 
    phi_stmt_2383_ack_6452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2383_ack_0, ack => convTransposeD_CP_5725_elements(83)); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_2297/merge_stmt_2382_PhiAck/phi_stmt_2389_ack
      -- 
    phi_stmt_2389_ack_6453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2389_ack_0, ack => convTransposeD_CP_5725_elements(84)); -- 
    -- CP-element group 85:  join  transition  place  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	89 
    -- CP-element group 85:  members (10) 
      -- CP-element group 85: 	 branch_block_stmt_2297/merge_stmt_2382__exit__
      -- CP-element group 85: 	 branch_block_stmt_2297/assign_stmt_2400_to_assign_stmt_2445__entry__
      -- CP-element group 85: 	 branch_block_stmt_2297/assign_stmt_2400_to_assign_stmt_2445__exit__
      -- CP-element group 85: 	 branch_block_stmt_2297/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 85: 	 branch_block_stmt_2297/assign_stmt_2400_to_assign_stmt_2445/$entry
      -- CP-element group 85: 	 branch_block_stmt_2297/assign_stmt_2400_to_assign_stmt_2445/$exit
      -- CP-element group 85: 	 branch_block_stmt_2297/merge_stmt_2382_PhiAck/$exit
      -- CP-element group 85: 	 branch_block_stmt_2297/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- CP-element group 85: 	 branch_block_stmt_2297/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2448/$entry
      -- CP-element group 85: 	 branch_block_stmt_2297/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/$entry
      -- 
    convTransposeD_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_5725_elements(83) & convTransposeD_CP_5725_elements(84);
      gj_convTransposeD_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_5725_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	56 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_2297/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/type_cast_2451/SplitProtocol/Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_2297/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/type_cast_2451/SplitProtocol/Sample/ra
      -- 
    ra_6473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2451_inst_ack_0, ack => convTransposeD_CP_5725_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	56 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_2297/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/type_cast_2451/SplitProtocol/Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_2297/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/type_cast_2451/SplitProtocol/Update/ca
      -- 
    ca_6478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2451_inst_ack_1, ack => convTransposeD_CP_5725_elements(87)); -- 
    -- CP-element group 88:  join  transition  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (6) 
      -- CP-element group 88: 	 branch_block_stmt_2297/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- CP-element group 88: 	 branch_block_stmt_2297/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2448/$exit
      -- CP-element group 88: 	 branch_block_stmt_2297/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/$exit
      -- CP-element group 88: 	 branch_block_stmt_2297/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/type_cast_2451/$exit
      -- CP-element group 88: 	 branch_block_stmt_2297/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/type_cast_2451/SplitProtocol/$exit
      -- CP-element group 88: 	 branch_block_stmt_2297/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2448/phi_stmt_2448_req
      -- 
    phi_stmt_2448_req_6479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2448_req_6479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(88), ack => phi_stmt_2448_req_0); -- 
    convTransposeD_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_5725_elements(86) & convTransposeD_CP_5725_elements(87);
      gj_convTransposeD_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_5725_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  transition  output  delay-element  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	85 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89:  members (5) 
      -- CP-element group 89: 	 branch_block_stmt_2297/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- CP-element group 89: 	 branch_block_stmt_2297/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2448/$exit
      -- CP-element group 89: 	 branch_block_stmt_2297/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/$exit
      -- CP-element group 89: 	 branch_block_stmt_2297/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/type_cast_2454_konst_delay_trans
      -- CP-element group 89: 	 branch_block_stmt_2297/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2448/phi_stmt_2448_req
      -- 
    phi_stmt_2448_req_6490_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2448_req_6490_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(89), ack => phi_stmt_2448_req_1); -- 
    -- Element group convTransposeD_CP_5725_elements(89) is a control-delay.
    cp_element_89_delay: control_delay_element  generic map(name => " 89_delay", delay_value => 1)  port map(req => convTransposeD_CP_5725_elements(85), ack => convTransposeD_CP_5725_elements(89), clk => clk, reset =>reset);
    -- CP-element group 90:  merge  transition  place  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_2297/merge_stmt_2447_PhiReqMerge
      -- CP-element group 90: 	 branch_block_stmt_2297/merge_stmt_2447_PhiAck/$entry
      -- 
    convTransposeD_CP_5725_elements(90) <= OrReduce(convTransposeD_CP_5725_elements(88) & convTransposeD_CP_5725_elements(89));
    -- CP-element group 91:  fork  transition  place  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	32 
    -- CP-element group 91: 	33 
    -- CP-element group 91: 	35 
    -- CP-element group 91: 	37 
    -- CP-element group 91: 	39 
    -- CP-element group 91: 	41 
    -- CP-element group 91: 	42 
    -- CP-element group 91: 	43 
    -- CP-element group 91: 	45 
    -- CP-element group 91: 	47 
    -- CP-element group 91: 	49 
    -- CP-element group 91: 	52 
    -- CP-element group 91: 	53 
    -- CP-element group 91: 	54 
    -- CP-element group 91:  members (51) 
      -- CP-element group 91: 	 branch_block_stmt_2297/merge_stmt_2447__exit__
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549__entry__
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/$entry
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2475_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2475_update_start_
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2475_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2475_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2475_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2475_Update/cr
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2489_update_start_
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2489_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2489_Update/cr
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/addr_of_2496_update_start_
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2495_final_index_sum_regn_update_start
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2495_final_index_sum_regn_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2495_final_index_sum_regn_Update/req
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/addr_of_2496_complete/$entry
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/addr_of_2496_complete/req
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2500_update_start_
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2500_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2500_Update/word_access_complete/$entry
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2500_Update/word_access_complete/word_0/$entry
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2500_Update/word_access_complete/word_0/cr
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2505_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2505_update_start_
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2505_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2505_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2505_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2505_Update/cr
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2519_update_start_
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2519_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2519_Update/cr
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/addr_of_2526_update_start_
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2525_final_index_sum_regn_update_start
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2525_final_index_sum_regn_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/array_obj_ref_2525_final_index_sum_regn_Update/req
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/addr_of_2526_complete/$entry
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/addr_of_2526_complete/req
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2529_update_start_
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2529_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2529_Update/word_access_complete/$entry
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2529_Update/word_access_complete/word_0/$entry
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/ptr_deref_2529_Update/word_access_complete/word_0/cr
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2535_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2535_update_start_
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2535_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2535_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2535_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_2297/assign_stmt_2461_to_assign_stmt_2549/type_cast_2535_Update/cr
      -- CP-element group 91: 	 branch_block_stmt_2297/merge_stmt_2447_PhiAck/$exit
      -- CP-element group 91: 	 branch_block_stmt_2297/merge_stmt_2447_PhiAck/phi_stmt_2448_ack
      -- 
    phi_stmt_2448_ack_6495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2448_ack_0, ack => convTransposeD_CP_5725_elements(91)); -- 
    rr_5992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(91), ack => type_cast_2475_inst_req_0); -- 
    cr_5997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(91), ack => type_cast_2475_inst_req_1); -- 
    cr_6011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(91), ack => type_cast_2489_inst_req_1); -- 
    req_6042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(91), ack => array_obj_ref_2495_index_offset_req_1); -- 
    req_6057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(91), ack => addr_of_2496_final_reg_req_1); -- 
    cr_6102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(91), ack => ptr_deref_2500_load_0_req_1); -- 
    rr_6116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(91), ack => type_cast_2505_inst_req_0); -- 
    cr_6121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(91), ack => type_cast_2505_inst_req_1); -- 
    cr_6135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(91), ack => type_cast_2519_inst_req_1); -- 
    req_6166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(91), ack => array_obj_ref_2525_index_offset_req_1); -- 
    req_6181_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6181_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(91), ack => addr_of_2526_final_reg_req_1); -- 
    cr_6231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(91), ack => ptr_deref_2529_store_0_req_1); -- 
    rr_6240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(91), ack => type_cast_2535_inst_req_0); -- 
    cr_6245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5725_elements(91), ack => type_cast_2535_inst_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_2483_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2513_wire : std_logic_vector(31 downto 0);
    signal R_idxprom102_2524_resized : std_logic_vector(13 downto 0);
    signal R_idxprom102_2524_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2494_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2494_scaled : std_logic_vector(13 downto 0);
    signal add107_2542 : std_logic_vector(31 downto 0);
    signal add49_2466 : std_logic_vector(15 downto 0);
    signal add93_2471 : std_logic_vector(15 downto 0);
    signal array_obj_ref_2495_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2495_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2495_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2495_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2495_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2495_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2525_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2525_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2525_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2525_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2525_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2525_root_address : std_logic_vector(13 downto 0);
    signal arrayidx103_2527 : std_logic_vector(31 downto 0);
    signal arrayidx97_2497 : std_logic_vector(31 downto 0);
    signal call11_2318 : std_logic_vector(15 downto 0);
    signal call13_2321 : std_logic_vector(15 downto 0);
    signal call14_2324 : std_logic_vector(15 downto 0);
    signal call15_2327 : std_logic_vector(15 downto 0);
    signal call17_2330 : std_logic_vector(15 downto 0);
    signal call19_2333 : std_logic_vector(15 downto 0);
    signal call1_2303 : std_logic_vector(15 downto 0);
    signal call3_2306 : std_logic_vector(15 downto 0);
    signal call5_2309 : std_logic_vector(15 downto 0);
    signal call7_2312 : std_logic_vector(15 downto 0);
    signal call9_2315 : std_logic_vector(15 downto 0);
    signal call_2300 : std_logic_vector(15 downto 0);
    signal cmp122_2580 : std_logic_vector(0 downto 0);
    signal cmp137_2605 : std_logic_vector(0 downto 0);
    signal cmp_2549 : std_logic_vector(0 downto 0);
    signal conv100_2506 : std_logic_vector(31 downto 0);
    signal conv106_2536 : std_logic_vector(31 downto 0);
    signal conv110_2350 : std_logic_vector(31 downto 0);
    signal conv118_2575 : std_logic_vector(31 downto 0);
    signal conv121_2354 : std_logic_vector(31 downto 0);
    signal conv133_2600 : std_logic_vector(31 downto 0);
    signal conv136_2358 : std_logic_vector(31 downto 0);
    signal conv96_2476 : std_logic_vector(31 downto 0);
    signal div27_2346 : std_logic_vector(15 downto 0);
    signal div_2340 : std_logic_vector(15 downto 0);
    signal idxprom102_2520 : std_logic_vector(63 downto 0);
    signal idxprom_2490 : std_logic_vector(63 downto 0);
    signal inc126_2590 : std_logic_vector(15 downto 0);
    signal inc_2570 : std_logic_vector(15 downto 0);
    signal indvar_2448 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_2562 : std_logic_vector(15 downto 0);
    signal input_dim0x_x0_2595 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_2389 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_2383 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2586 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2461 : std_logic_vector(15 downto 0);
    signal ptr_deref_2500_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2500_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2500_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2500_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2500_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2529_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2529_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2529_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2529_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2529_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2529_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr101_2515 : std_logic_vector(31 downto 0);
    signal shr_2485 : std_logic_vector(31 downto 0);
    signal tmp10_2445 : std_logic_vector(15 downto 0);
    signal tmp164_2400 : std_logic_vector(15 downto 0);
    signal tmp165_2405 : std_logic_vector(15 downto 0);
    signal tmp166_2410 : std_logic_vector(15 downto 0);
    signal tmp1_2369 : std_logic_vector(15 downto 0);
    signal tmp2_2415 : std_logic_vector(15 downto 0);
    signal tmp3_2420 : std_logic_vector(15 downto 0);
    signal tmp4_2375 : std_logic_vector(15 downto 0);
    signal tmp5_2380 : std_logic_vector(15 downto 0);
    signal tmp6_2425 : std_logic_vector(15 downto 0);
    signal tmp7_2430 : std_logic_vector(15 downto 0);
    signal tmp8_2435 : std_logic_vector(15 downto 0);
    signal tmp98_2501 : std_logic_vector(63 downto 0);
    signal tmp9_2440 : std_logic_vector(15 downto 0);
    signal tmp_2364 : std_logic_vector(15 downto 0);
    signal type_cast_2338_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2344_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2362_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2373_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2386_wire : std_logic_vector(15 downto 0);
    signal type_cast_2388_wire : std_logic_vector(15 downto 0);
    signal type_cast_2392_wire : std_logic_vector(15 downto 0);
    signal type_cast_2394_wire : std_logic_vector(15 downto 0);
    signal type_cast_2451_wire : std_logic_vector(15 downto 0);
    signal type_cast_2454_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2459_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2474_wire : std_logic_vector(31 downto 0);
    signal type_cast_2479_wire : std_logic_vector(31 downto 0);
    signal type_cast_2482_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2488_wire : std_logic_vector(63 downto 0);
    signal type_cast_2504_wire : std_logic_vector(31 downto 0);
    signal type_cast_2509_wire : std_logic_vector(31 downto 0);
    signal type_cast_2512_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2518_wire : std_logic_vector(63 downto 0);
    signal type_cast_2534_wire : std_logic_vector(31 downto 0);
    signal type_cast_2540_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2545_wire : std_logic_vector(31 downto 0);
    signal type_cast_2547_wire : std_logic_vector(31 downto 0);
    signal type_cast_2560_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2568_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2573_wire : std_logic_vector(31 downto 0);
    signal type_cast_2598_wire : std_logic_vector(31 downto 0);
    signal type_cast_2616_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_2495_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2495_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2495_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2495_resized_base_address <= "00000000000000";
    array_obj_ref_2525_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2525_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2525_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2525_resized_base_address <= "00000000000000";
    ptr_deref_2500_word_offset_0 <= "00000000000000";
    ptr_deref_2529_word_offset_0 <= "00000000000000";
    type_cast_2338_wire_constant <= "0000000000000001";
    type_cast_2344_wire_constant <= "0000000000000001";
    type_cast_2362_wire_constant <= "1111111111111111";
    type_cast_2373_wire_constant <= "1111111111111111";
    type_cast_2454_wire_constant <= "0000000000000000";
    type_cast_2459_wire_constant <= "0000000000000100";
    type_cast_2482_wire_constant <= "00000000000000000000000000000010";
    type_cast_2512_wire_constant <= "00000000000000000000000000000010";
    type_cast_2540_wire_constant <= "00000000000000000000000000000100";
    type_cast_2560_wire_constant <= "0000000000000001";
    type_cast_2568_wire_constant <= "0000000000000001";
    type_cast_2616_wire_constant <= "0000000000000001";
    phi_stmt_2383: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2386_wire & type_cast_2388_wire;
      req <= phi_stmt_2383_req_0 & phi_stmt_2383_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2383",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2383_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_2383,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2383
    phi_stmt_2389: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2392_wire & type_cast_2394_wire;
      req <= phi_stmt_2389_req_0 & phi_stmt_2389_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2389",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2389_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_2389,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2389
    phi_stmt_2448: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2451_wire & type_cast_2454_wire_constant;
      req <= phi_stmt_2448_req_0 & phi_stmt_2448_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2448",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2448_ack_0,
          idata => idata,
          odata => indvar_2448,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2448
    -- flow-through select operator MUX_2585_inst
    input_dim1x_x2_2586 <= div27_2346 when (cmp122_2580(0) /=  '0') else inc_2570;
    addr_of_2496_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2496_final_reg_req_0;
      addr_of_2496_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2496_final_reg_req_1;
      addr_of_2496_final_reg_ack_1<= rack(0);
      addr_of_2496_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2496_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2495_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx97_2497,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2526_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2526_final_reg_req_0;
      addr_of_2526_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2526_final_reg_req_1;
      addr_of_2526_final_reg_ack_1<= rack(0);
      addr_of_2526_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2526_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2525_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx103_2527,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2349_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2349_inst_req_0;
      type_cast_2349_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2349_inst_req_1;
      type_cast_2349_inst_ack_1<= rack(0);
      type_cast_2349_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2349_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_2306,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv110_2350,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2353_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2353_inst_req_0;
      type_cast_2353_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2353_inst_req_1;
      type_cast_2353_inst_ack_1<= rack(0);
      type_cast_2353_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2353_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1_2303,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv121_2354,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2357_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2357_inst_req_0;
      type_cast_2357_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2357_inst_req_1;
      type_cast_2357_inst_ack_1<= rack(0);
      type_cast_2357_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2357_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_2300,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv136_2358,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2386_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2386_inst_req_0;
      type_cast_2386_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2386_inst_req_1;
      type_cast_2386_inst_ack_1<= rack(0);
      type_cast_2386_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2386_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div27_2346,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2386_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2388_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2388_inst_req_0;
      type_cast_2388_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2388_inst_req_1;
      type_cast_2388_inst_ack_1<= rack(0);
      type_cast_2388_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2388_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2586,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2388_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2392_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2392_inst_req_0;
      type_cast_2392_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2392_inst_req_1;
      type_cast_2392_inst_ack_1<= rack(0);
      type_cast_2392_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2392_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x0_2595,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2392_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2394_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2394_inst_req_0;
      type_cast_2394_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2394_inst_req_1;
      type_cast_2394_inst_ack_1<= rack(0);
      type_cast_2394_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2394_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_2340,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2394_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2451_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2451_inst_req_0;
      type_cast_2451_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2451_inst_req_1;
      type_cast_2451_inst_ack_1<= rack(0);
      type_cast_2451_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2451_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2562,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2451_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2475_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2475_inst_req_0;
      type_cast_2475_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2475_inst_req_1;
      type_cast_2475_inst_ack_1<= rack(0);
      type_cast_2475_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2475_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2474_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv96_2476,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2479_inst
    process(conv96_2476) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv96_2476(31 downto 0);
      type_cast_2479_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2484_inst
    process(ASHR_i32_i32_2483_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2483_wire(31 downto 0);
      shr_2485 <= tmp_var; -- 
    end process;
    type_cast_2489_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2489_inst_req_0;
      type_cast_2489_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2489_inst_req_1;
      type_cast_2489_inst_ack_1<= rack(0);
      type_cast_2489_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2489_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2488_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2490,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2505_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2505_inst_req_0;
      type_cast_2505_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2505_inst_req_1;
      type_cast_2505_inst_ack_1<= rack(0);
      type_cast_2505_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2505_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2504_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv100_2506,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2509_inst
    process(conv100_2506) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv100_2506(31 downto 0);
      type_cast_2509_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2514_inst
    process(ASHR_i32_i32_2513_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2513_wire(31 downto 0);
      shr101_2515 <= tmp_var; -- 
    end process;
    type_cast_2519_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2519_inst_req_0;
      type_cast_2519_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2519_inst_req_1;
      type_cast_2519_inst_ack_1<= rack(0);
      type_cast_2519_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2519_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2518_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom102_2520,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2535_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2535_inst_req_0;
      type_cast_2535_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2535_inst_req_1;
      type_cast_2535_inst_ack_1<= rack(0);
      type_cast_2535_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2535_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2534_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv106_2536,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2545_inst
    process(add107_2542) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add107_2542(31 downto 0);
      type_cast_2545_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2547_inst
    process(conv110_2350) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv110_2350(31 downto 0);
      type_cast_2547_wire <= tmp_var; -- 
    end process;
    type_cast_2574_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2574_inst_req_0;
      type_cast_2574_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2574_inst_req_1;
      type_cast_2574_inst_ack_1<= rack(0);
      type_cast_2574_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2574_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2573_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv118_2575,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2589_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2589_inst_req_0;
      type_cast_2589_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2589_inst_req_1;
      type_cast_2589_inst_ack_1<= rack(0);
      type_cast_2589_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2589_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp122_2580,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc126_2590,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2599_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2599_inst_req_0;
      type_cast_2599_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2599_inst_req_1;
      type_cast_2599_inst_ack_1<= rack(0);
      type_cast_2599_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2599_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2598_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv133_2600,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_2495_index_1_rename
    process(R_idxprom_2494_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2494_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2494_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2495_index_1_resize
    process(idxprom_2490) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2490;
      ov := iv(13 downto 0);
      R_idxprom_2494_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2495_root_address_inst
    process(array_obj_ref_2495_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2495_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2495_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2525_index_1_rename
    process(R_idxprom102_2524_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom102_2524_resized;
      ov(13 downto 0) := iv;
      R_idxprom102_2524_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2525_index_1_resize
    process(idxprom102_2520) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom102_2520;
      ov := iv(13 downto 0);
      R_idxprom102_2524_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2525_root_address_inst
    process(array_obj_ref_2525_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2525_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2525_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2500_addr_0
    process(ptr_deref_2500_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2500_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2500_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2500_base_resize
    process(arrayidx97_2497) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx97_2497;
      ov := iv(13 downto 0);
      ptr_deref_2500_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2500_gather_scatter
    process(ptr_deref_2500_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2500_data_0;
      ov(63 downto 0) := iv;
      tmp98_2501 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2500_root_address_inst
    process(ptr_deref_2500_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2500_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2500_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2529_addr_0
    process(ptr_deref_2529_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2529_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2529_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2529_base_resize
    process(arrayidx103_2527) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx103_2527;
      ov := iv(13 downto 0);
      ptr_deref_2529_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2529_gather_scatter
    process(tmp98_2501) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp98_2501;
      ov(63 downto 0) := iv;
      ptr_deref_2529_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2529_root_address_inst
    process(ptr_deref_2529_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2529_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2529_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2550_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2549;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2550_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2550_branch_req_0,
          ack0 => if_stmt_2550_branch_ack_0,
          ack1 => if_stmt_2550_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2606_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp137_2605;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2606_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2606_branch_req_0,
          ack0 => if_stmt_2606_branch_ack_0,
          ack1 => if_stmt_2606_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2363_inst
    process(call9_2315) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_2315, type_cast_2362_wire_constant, tmp_var);
      tmp_2364 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2374_inst
    process(call7_2312) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_2312, type_cast_2373_wire_constant, tmp_var);
      tmp4_2375 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2404_inst
    process(input_dim1x_x1x_xph_2383, tmp164_2400) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_2383, tmp164_2400, tmp_var);
      tmp165_2405 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2419_inst
    process(tmp1_2369, tmp2_2415) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp1_2369, tmp2_2415, tmp_var);
      tmp3_2420 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2429_inst
    process(tmp5_2380, tmp6_2425) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp5_2380, tmp6_2425, tmp_var);
      tmp7_2430 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2439_inst
    process(tmp3_2420, tmp8_2435) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp3_2420, tmp8_2435, tmp_var);
      tmp9_2440 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2465_inst
    process(tmp166_2410, input_dim2x_x1_2461) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp166_2410, input_dim2x_x1_2461, tmp_var);
      add49_2466 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2470_inst
    process(tmp10_2445, input_dim2x_x1_2461) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp10_2445, input_dim2x_x1_2461, tmp_var);
      add93_2471 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2561_inst
    process(indvar_2448) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2448, type_cast_2560_wire_constant, tmp_var);
      indvarx_xnext_2562 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2569_inst
    process(input_dim1x_x1x_xph_2383) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_2383, type_cast_2568_wire_constant, tmp_var);
      inc_2570 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2594_inst
    process(inc126_2590, input_dim0x_x2x_xph_2389) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc126_2590, input_dim0x_x2x_xph_2389, tmp_var);
      input_dim0x_x0_2595 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2541_inst
    process(conv106_2536) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv106_2536, type_cast_2540_wire_constant, tmp_var);
      add107_2542 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2483_inst
    process(type_cast_2479_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2479_wire, type_cast_2482_wire_constant, tmp_var);
      ASHR_i32_i32_2483_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2513_inst
    process(type_cast_2509_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2509_wire, type_cast_2512_wire_constant, tmp_var);
      ASHR_i32_i32_2513_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2579_inst
    process(conv118_2575, conv121_2354) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv118_2575, conv121_2354, tmp_var);
      cmp122_2580 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2604_inst
    process(conv133_2600, conv136_2358) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv133_2600, conv136_2358, tmp_var);
      cmp137_2605 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2339_inst
    process(call_2300) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_2300, type_cast_2338_wire_constant, tmp_var);
      div_2340 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2345_inst
    process(call1_2303) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call1_2303, type_cast_2344_wire_constant, tmp_var);
      div27_2346 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2399_inst
    process(call1_2303, input_dim0x_x2x_xph_2389) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call1_2303, input_dim0x_x2x_xph_2389, tmp_var);
      tmp164_2400 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2409_inst
    process(call3_2306, tmp165_2405) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call3_2306, tmp165_2405, tmp_var);
      tmp166_2410 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2414_inst
    process(call13_2321, input_dim1x_x1x_xph_2383) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call13_2321, input_dim1x_x1x_xph_2383, tmp_var);
      tmp2_2415 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2424_inst
    process(call13_2321, input_dim0x_x2x_xph_2389) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call13_2321, input_dim0x_x2x_xph_2389, tmp_var);
      tmp6_2425 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2434_inst
    process(call17_2330, tmp7_2430) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call17_2330, tmp7_2430, tmp_var);
      tmp8_2435 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2444_inst
    process(call19_2333, tmp9_2440) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call19_2333, tmp9_2440, tmp_var);
      tmp10_2445 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2460_inst
    process(indvar_2448) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2448, type_cast_2459_wire_constant, tmp_var);
      input_dim2x_x1_2461 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2548_inst
    process(type_cast_2545_wire, type_cast_2547_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2545_wire, type_cast_2547_wire, tmp_var);
      cmp_2549 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2368_inst
    process(tmp_2364, call14_2324) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp_2364, call14_2324, tmp_var);
      tmp1_2369 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2379_inst
    process(tmp4_2375, call14_2324) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp4_2375, call14_2324, tmp_var);
      tmp5_2380 <= tmp_var; --
    end process;
    -- shared split operator group (28) : array_obj_ref_2495_index_offset 
    ApIntAdd_group_28: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2494_scaled;
      array_obj_ref_2495_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2495_index_offset_req_0;
      array_obj_ref_2495_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2495_index_offset_req_1;
      array_obj_ref_2495_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_28_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_28_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : array_obj_ref_2525_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom102_2524_scaled;
      array_obj_ref_2525_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2525_index_offset_req_0;
      array_obj_ref_2525_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2525_index_offset_req_1;
      array_obj_ref_2525_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- unary operator type_cast_2474_inst
    process(add49_2466) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", add49_2466, tmp_var);
      type_cast_2474_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2488_inst
    process(shr_2485) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_2485, tmp_var);
      type_cast_2488_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2504_inst
    process(add93_2471) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", add93_2471, tmp_var);
      type_cast_2504_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2518_inst
    process(shr101_2515) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr101_2515, tmp_var);
      type_cast_2518_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2534_inst
    process(input_dim2x_x1_2461) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim2x_x1_2461, tmp_var);
      type_cast_2534_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2573_inst
    process(inc_2570) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_2570, tmp_var);
      type_cast_2573_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2598_inst
    process(input_dim0x_x0_2595) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim0x_x0_2595, tmp_var);
      type_cast_2598_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_2500_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2500_load_0_req_0;
      ptr_deref_2500_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2500_load_0_req_1;
      ptr_deref_2500_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2500_word_address_0;
      ptr_deref_2500_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_2529_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2529_store_0_req_0;
      ptr_deref_2529_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2529_store_0_req_1;
      ptr_deref_2529_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2529_word_address_0;
      data_in <= ptr_deref_2529_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block1_start_2323_inst RPIPE_Block1_start_2326_inst RPIPE_Block1_start_2329_inst RPIPE_Block1_start_2332_inst RPIPE_Block1_start_2320_inst RPIPE_Block1_start_2317_inst RPIPE_Block1_start_2314_inst RPIPE_Block1_start_2311_inst RPIPE_Block1_start_2308_inst RPIPE_Block1_start_2305_inst RPIPE_Block1_start_2302_inst RPIPE_Block1_start_2299_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(191 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 11 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 11 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 11 downto 0);
      signal guard_vector : std_logic_vector( 11 downto 0);
      constant outBUFs : IntegerArray(11 downto 0) := (11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(11 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false);
      constant guardBuffering: IntegerArray(11 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2);
      -- 
    begin -- 
      reqL_unguarded(11) <= RPIPE_Block1_start_2323_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block1_start_2326_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block1_start_2329_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block1_start_2332_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block1_start_2320_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block1_start_2317_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block1_start_2314_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block1_start_2311_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block1_start_2308_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block1_start_2305_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block1_start_2302_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block1_start_2299_inst_req_0;
      RPIPE_Block1_start_2323_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block1_start_2326_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block1_start_2329_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block1_start_2332_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block1_start_2320_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block1_start_2317_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block1_start_2314_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block1_start_2311_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block1_start_2308_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block1_start_2305_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block1_start_2302_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block1_start_2299_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(11) <= RPIPE_Block1_start_2323_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block1_start_2326_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block1_start_2329_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block1_start_2332_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block1_start_2320_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block1_start_2317_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block1_start_2314_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block1_start_2311_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block1_start_2308_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block1_start_2305_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block1_start_2302_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block1_start_2299_inst_req_1;
      RPIPE_Block1_start_2323_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block1_start_2326_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block1_start_2329_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block1_start_2332_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block1_start_2320_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block1_start_2317_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block1_start_2314_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block1_start_2311_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block1_start_2308_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block1_start_2305_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block1_start_2302_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block1_start_2299_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      call14_2324 <= data_out(191 downto 176);
      call15_2327 <= data_out(175 downto 160);
      call17_2330 <= data_out(159 downto 144);
      call19_2333 <= data_out(143 downto 128);
      call13_2321 <= data_out(127 downto 112);
      call11_2318 <= data_out(111 downto 96);
      call9_2315 <= data_out(95 downto 80);
      call7_2312 <= data_out(79 downto 64);
      call5_2309 <= data_out(63 downto 48);
      call3_2306 <= data_out(47 downto 32);
      call1_2303 <= data_out(31 downto 16);
      call_2300 <= data_out(15 downto 0);
      Block1_start_read_0_gI: SplitGuardInterface generic map(name => "Block1_start_read_0_gI", nreqs => 12, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_start_read_0: InputPortRevised -- 
        generic map ( name => "Block1_start_read_0", data_width => 16,  num_reqs => 12,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_start_pipe_read_req(0),
          oack => Block1_start_pipe_read_ack(0),
          odata => Block1_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block3_done_2614_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block3_done_2614_inst_req_0;
      WPIPE_Block3_done_2614_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block3_done_2614_inst_req_1;
      WPIPE_Block3_done_2614_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2616_wire_constant;
      Block3_done_write_0_gI: SplitGuardInterface generic map(name => "Block3_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block3_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_done_pipe_write_req(0),
          oack => Block3_done_pipe_write_ack(0),
          odata => Block3_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeD_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    c : out  std_logic_vector(63 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal c_buffer :  std_logic_vector(63 downto 0);
  signal c_update_enable: Boolean;
  signal timer_CP_0_start: Boolean;
  signal timer_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal LOAD_count_29_load_0_req_0 : boolean;
  signal LOAD_count_29_load_0_ack_0 : boolean;
  signal LOAD_count_29_load_0_req_1 : boolean;
  signal LOAD_count_29_load_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= c_buffer;
  c <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_0: Block -- control-path 
    signal timer_CP_0_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    timer_CP_0_elements(0) <= timer_CP_0_start;
    timer_CP_0_symbol <= timer_CP_0_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_Update/$entry
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_30/$entry
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_sample_start_
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_update_start_
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_Sample/$entry
      -- 
    cr_32_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_32_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => LOAD_count_29_load_0_req_1); -- 
    rr_21_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_21_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => LOAD_count_29_load_0_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 assign_stmt_30/LOAD_count_29_Sample/word_access_start/$exit
      -- CP-element group 1: 	 assign_stmt_30/LOAD_count_29_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 assign_stmt_30/LOAD_count_29_Sample/word_access_start/word_0/ra
      -- CP-element group 1: 	 assign_stmt_30/LOAD_count_29_sample_completed_
      -- CP-element group 1: 	 assign_stmt_30/LOAD_count_29_Sample/$exit
      -- 
    ra_22_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_29_load_0_ack_0, ack => timer_CP_0_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_Update/$exit
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_Update/word_access_complete/$exit
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_Update/LOAD_count_29_Merge/$entry
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_30/$exit
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_update_completed_
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_Update/LOAD_count_29_Merge/$exit
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_Update/LOAD_count_29_Merge/merge_req
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_Update/LOAD_count_29_Merge/merge_ack
      -- 
    ca_33_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_29_load_0_ack_1, ack => timer_CP_0_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_count_29_data_0 : std_logic_vector(63 downto 0);
    signal LOAD_count_29_word_address_0 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    LOAD_count_29_word_address_0 <= "0";
    -- equivalence LOAD_count_29_gather_scatter
    process(LOAD_count_29_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_count_29_data_0;
      ov(63 downto 0) := iv;
      c_buffer <= ov(63 downto 0);
      --
    end process;
    -- shared load operator group (0) : LOAD_count_29_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_count_29_load_0_req_0;
      LOAD_count_29_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_count_29_load_0_req_1;
      LOAD_count_29_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_count_29_word_address_0;
      LOAD_count_29_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(0 downto 0),
          mtag => memory_space_0_lr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    Block2_start_pipe_read_data: out std_logic_vector(15 downto 0);
    Block2_start_pipe_read_req : in std_logic_vector(0 downto 0);
    Block2_start_pipe_read_ack : out std_logic_vector(0 downto 0);
    Block3_start_pipe_read_data: out std_logic_vector(15 downto 0);
    Block3_start_pipe_read_req : in std_logic_vector(0 downto 0);
    Block3_start_pipe_read_ack : out std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    ConvTranspose_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    ConvTranspose_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_read_data: out std_logic_vector(63 downto 0);
    elapsed_time_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(55 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(75 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(255 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(10 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_3
  signal memory_space_3_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_3_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_3_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_3_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_3_sr_req :  std_logic_vector(4 downto 0);
  signal memory_space_3_sr_ack : std_logic_vector(4 downto 0);
  signal memory_space_3_sr_addr : std_logic_vector(69 downto 0);
  signal memory_space_3_sr_data : std_logic_vector(319 downto 0);
  signal memory_space_3_sr_tag : std_logic_vector(94 downto 0);
  signal memory_space_3_sc_req : std_logic_vector(4 downto 0);
  signal memory_space_3_sc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_3_sc_tag :  std_logic_vector(4 downto 0);
  -- declarations related to module convTranspose
  component convTranspose is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTranspose
  signal convTranspose_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTranspose_tag_out   : std_logic_vector(1 downto 0);
  signal convTranspose_start_req : std_logic;
  signal convTranspose_start_ack : std_logic;
  signal convTranspose_fin_req   : std_logic;
  signal convTranspose_fin_ack : std_logic;
  -- declarations related to module convTransposeA
  component convTransposeA is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeA
  signal convTransposeA_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeA_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeA_start_req : std_logic;
  signal convTransposeA_start_ack : std_logic;
  signal convTransposeA_fin_req   : std_logic;
  signal convTransposeA_fin_ack : std_logic;
  -- declarations related to module convTransposeB
  component convTransposeB is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeB
  signal convTransposeB_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeB_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeB_start_req : std_logic;
  signal convTransposeB_start_ack : std_logic;
  signal convTransposeB_fin_req   : std_logic;
  signal convTransposeB_fin_ack : std_logic;
  -- declarations related to module convTransposeC
  component convTransposeC is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeC
  signal convTransposeC_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeC_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeC_start_req : std_logic;
  signal convTransposeC_start_ack : std_logic;
  signal convTransposeC_fin_req   : std_logic;
  signal convTransposeC_fin_ack : std_logic;
  -- declarations related to module convTransposeD
  component convTransposeD is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeD
  signal convTransposeD_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeD_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeD_start_req : std_logic;
  signal convTransposeD_start_ack : std_logic;
  signal convTransposeD_fin_req   : std_logic;
  signal convTransposeD_fin_ack : std_logic;
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_c :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe Block0_done
  signal Block0_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_done
  signal Block0_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block0_start
  signal Block0_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_start
  signal Block0_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_done
  signal Block1_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_done
  signal Block1_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_start
  signal Block1_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_start
  signal Block1_start_pipe_read_data: std_logic_vector(47 downto 0);
  signal Block1_start_pipe_read_req: std_logic_vector(2 downto 0);
  signal Block1_start_pipe_read_ack: std_logic_vector(2 downto 0);
  -- aggregate signals for write to pipe Block2_done
  signal Block2_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_done
  signal Block2_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_start
  signal Block2_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_done
  signal Block3_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_done
  signal Block3_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_start
  signal Block3_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe ConvTranspose_input_pipe
  signal ConvTranspose_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe ConvTranspose_output_pipe
  signal ConvTranspose_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe elapsed_time_pipe
  signal elapsed_time_pipe_pipe_write_data: std_logic_vector(63 downto 0);
  signal elapsed_time_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal elapsed_time_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module convTranspose
  convTranspose_instance:convTranspose-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTranspose_start_req,
      start_ack => convTranspose_start_ack,
      fin_req => convTranspose_fin_req,
      fin_ack => convTranspose_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_3_lr_req => memory_space_3_lr_req(0 downto 0),
      memory_space_3_lr_ack => memory_space_3_lr_ack(0 downto 0),
      memory_space_3_lr_addr => memory_space_3_lr_addr(13 downto 0),
      memory_space_3_lr_tag => memory_space_3_lr_tag(18 downto 0),
      memory_space_3_lc_req => memory_space_3_lc_req(0 downto 0),
      memory_space_3_lc_ack => memory_space_3_lc_ack(0 downto 0),
      memory_space_3_lc_data => memory_space_3_lc_data(63 downto 0),
      memory_space_3_lc_tag => memory_space_3_lc_tag(0 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(18 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(0 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(10 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(63 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(0 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(0 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(4 downto 4),
      memory_space_3_sr_ack => memory_space_3_sr_ack(4 downto 4),
      memory_space_3_sr_addr => memory_space_3_sr_addr(69 downto 56),
      memory_space_3_sr_data => memory_space_3_sr_data(319 downto 256),
      memory_space_3_sr_tag => memory_space_3_sr_tag(94 downto 76),
      memory_space_3_sc_req => memory_space_3_sc_req(4 downto 4),
      memory_space_3_sc_ack => memory_space_3_sc_ack(4 downto 4),
      memory_space_3_sc_tag => memory_space_3_sc_tag(4 downto 4),
      Block0_done_pipe_read_req => Block0_done_pipe_read_req(0 downto 0),
      Block0_done_pipe_read_ack => Block0_done_pipe_read_ack(0 downto 0),
      Block0_done_pipe_read_data => Block0_done_pipe_read_data(15 downto 0),
      Block1_done_pipe_read_req => Block1_done_pipe_read_req(0 downto 0),
      Block1_done_pipe_read_ack => Block1_done_pipe_read_ack(0 downto 0),
      Block1_done_pipe_read_data => Block1_done_pipe_read_data(15 downto 0),
      ConvTranspose_input_pipe_pipe_read_req => ConvTranspose_input_pipe_pipe_read_req(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_ack => ConvTranspose_input_pipe_pipe_read_ack(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_data => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
      Block2_done_pipe_read_req => Block2_done_pipe_read_req(0 downto 0),
      Block2_done_pipe_read_ack => Block2_done_pipe_read_ack(0 downto 0),
      Block2_done_pipe_read_data => Block2_done_pipe_read_data(15 downto 0),
      Block3_done_pipe_read_req => Block3_done_pipe_read_req(0 downto 0),
      Block3_done_pipe_read_ack => Block3_done_pipe_read_ack(0 downto 0),
      Block3_done_pipe_read_data => Block3_done_pipe_read_data(15 downto 0),
      Block1_start_pipe_write_req => Block1_start_pipe_write_req(0 downto 0),
      Block1_start_pipe_write_ack => Block1_start_pipe_write_ack(0 downto 0),
      Block1_start_pipe_write_data => Block1_start_pipe_write_data(15 downto 0),
      Block0_start_pipe_write_req => Block0_start_pipe_write_req(0 downto 0),
      Block0_start_pipe_write_ack => Block0_start_pipe_write_ack(0 downto 0),
      Block0_start_pipe_write_data => Block0_start_pipe_write_data(15 downto 0),
      Block3_start_pipe_write_req => Block3_start_pipe_write_req(0 downto 0),
      Block3_start_pipe_write_ack => Block3_start_pipe_write_ack(0 downto 0),
      Block3_start_pipe_write_data => Block3_start_pipe_write_data(15 downto 0),
      ConvTranspose_output_pipe_pipe_write_req => ConvTranspose_output_pipe_pipe_write_req(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_ack => ConvTranspose_output_pipe_pipe_write_ack(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_data => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
      Block2_start_pipe_write_req => Block2_start_pipe_write_req(0 downto 0),
      Block2_start_pipe_write_ack => Block2_start_pipe_write_ack(0 downto 0),
      Block2_start_pipe_write_data => Block2_start_pipe_write_data(15 downto 0),
      elapsed_time_pipe_pipe_write_req => elapsed_time_pipe_pipe_write_req(0 downto 0),
      elapsed_time_pipe_pipe_write_ack => elapsed_time_pipe_pipe_write_ack(0 downto 0),
      elapsed_time_pipe_pipe_write_data => elapsed_time_pipe_pipe_write_data(63 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      tag_in => convTranspose_tag_in,
      tag_out => convTranspose_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTranspose_tag_in <= (others => '0');
  convTranspose_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTranspose_start_req, start_ack => convTranspose_start_ack,  fin_req => convTranspose_fin_req,  fin_ack => convTranspose_fin_ack);
  -- module convTransposeA
  convTransposeA_instance:convTransposeA-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeA_start_req,
      start_ack => convTransposeA_start_ack,
      fin_req => convTransposeA_fin_req,
      fin_ack => convTransposeA_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(3 downto 3),
      memory_space_1_lr_ack => memory_space_1_lr_ack(3 downto 3),
      memory_space_1_lr_addr => memory_space_1_lr_addr(55 downto 42),
      memory_space_1_lr_tag => memory_space_1_lr_tag(75 downto 57),
      memory_space_1_lc_req => memory_space_1_lc_req(3 downto 3),
      memory_space_1_lc_ack => memory_space_1_lc_ack(3 downto 3),
      memory_space_1_lc_data => memory_space_1_lc_data(255 downto 192),
      memory_space_1_lc_tag => memory_space_1_lc_tag(3 downto 3),
      memory_space_3_sr_req => memory_space_3_sr_req(3 downto 3),
      memory_space_3_sr_ack => memory_space_3_sr_ack(3 downto 3),
      memory_space_3_sr_addr => memory_space_3_sr_addr(55 downto 42),
      memory_space_3_sr_data => memory_space_3_sr_data(255 downto 192),
      memory_space_3_sr_tag => memory_space_3_sr_tag(75 downto 57),
      memory_space_3_sc_req => memory_space_3_sc_req(3 downto 3),
      memory_space_3_sc_ack => memory_space_3_sc_ack(3 downto 3),
      memory_space_3_sc_tag => memory_space_3_sc_tag(3 downto 3),
      Block0_start_pipe_read_req => Block0_start_pipe_read_req(0 downto 0),
      Block0_start_pipe_read_ack => Block0_start_pipe_read_ack(0 downto 0),
      Block0_start_pipe_read_data => Block0_start_pipe_read_data(15 downto 0),
      Block0_done_pipe_write_req => Block0_done_pipe_write_req(0 downto 0),
      Block0_done_pipe_write_ack => Block0_done_pipe_write_ack(0 downto 0),
      Block0_done_pipe_write_data => Block0_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeA_tag_in,
      tag_out => convTransposeA_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeA_tag_in <= (others => '0');
  convTransposeA_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeA_start_req, start_ack => convTransposeA_start_ack,  fin_req => convTransposeA_fin_req,  fin_ack => convTransposeA_fin_ack);
  -- module convTransposeB
  convTransposeB_instance:convTransposeB-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeB_start_req,
      start_ack => convTransposeB_start_ack,
      fin_req => convTransposeB_fin_req,
      fin_ack => convTransposeB_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(1 downto 1),
      memory_space_1_lr_ack => memory_space_1_lr_ack(1 downto 1),
      memory_space_1_lr_addr => memory_space_1_lr_addr(27 downto 14),
      memory_space_1_lr_tag => memory_space_1_lr_tag(37 downto 19),
      memory_space_1_lc_req => memory_space_1_lc_req(1 downto 1),
      memory_space_1_lc_ack => memory_space_1_lc_ack(1 downto 1),
      memory_space_1_lc_data => memory_space_1_lc_data(127 downto 64),
      memory_space_1_lc_tag => memory_space_1_lc_tag(1 downto 1),
      memory_space_3_sr_req => memory_space_3_sr_req(1 downto 1),
      memory_space_3_sr_ack => memory_space_3_sr_ack(1 downto 1),
      memory_space_3_sr_addr => memory_space_3_sr_addr(27 downto 14),
      memory_space_3_sr_data => memory_space_3_sr_data(127 downto 64),
      memory_space_3_sr_tag => memory_space_3_sr_tag(37 downto 19),
      memory_space_3_sc_req => memory_space_3_sc_req(1 downto 1),
      memory_space_3_sc_ack => memory_space_3_sc_ack(1 downto 1),
      memory_space_3_sc_tag => memory_space_3_sc_tag(1 downto 1),
      Block1_start_pipe_read_req => Block1_start_pipe_read_req(1 downto 1),
      Block1_start_pipe_read_ack => Block1_start_pipe_read_ack(1 downto 1),
      Block1_start_pipe_read_data => Block1_start_pipe_read_data(31 downto 16),
      Block1_done_pipe_write_req => Block1_done_pipe_write_req(0 downto 0),
      Block1_done_pipe_write_ack => Block1_done_pipe_write_ack(0 downto 0),
      Block1_done_pipe_write_data => Block1_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeB_tag_in,
      tag_out => convTransposeB_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeB_tag_in <= (others => '0');
  convTransposeB_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeB_start_req, start_ack => convTransposeB_start_ack,  fin_req => convTransposeB_fin_req,  fin_ack => convTransposeB_fin_ack);
  -- module convTransposeC
  convTransposeC_instance:convTransposeC-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeC_start_req,
      start_ack => convTransposeC_start_ack,
      fin_req => convTransposeC_fin_req,
      fin_ack => convTransposeC_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(2 downto 2),
      memory_space_1_lr_ack => memory_space_1_lr_ack(2 downto 2),
      memory_space_1_lr_addr => memory_space_1_lr_addr(41 downto 28),
      memory_space_1_lr_tag => memory_space_1_lr_tag(56 downto 38),
      memory_space_1_lc_req => memory_space_1_lc_req(2 downto 2),
      memory_space_1_lc_ack => memory_space_1_lc_ack(2 downto 2),
      memory_space_1_lc_data => memory_space_1_lc_data(191 downto 128),
      memory_space_1_lc_tag => memory_space_1_lc_tag(2 downto 2),
      memory_space_3_sr_req => memory_space_3_sr_req(2 downto 2),
      memory_space_3_sr_ack => memory_space_3_sr_ack(2 downto 2),
      memory_space_3_sr_addr => memory_space_3_sr_addr(41 downto 28),
      memory_space_3_sr_data => memory_space_3_sr_data(191 downto 128),
      memory_space_3_sr_tag => memory_space_3_sr_tag(56 downto 38),
      memory_space_3_sc_req => memory_space_3_sc_req(2 downto 2),
      memory_space_3_sc_ack => memory_space_3_sc_ack(2 downto 2),
      memory_space_3_sc_tag => memory_space_3_sc_tag(2 downto 2),
      Block1_start_pipe_read_req => Block1_start_pipe_read_req(2 downto 2),
      Block1_start_pipe_read_ack => Block1_start_pipe_read_ack(2 downto 2),
      Block1_start_pipe_read_data => Block1_start_pipe_read_data(47 downto 32),
      Block2_done_pipe_write_req => Block2_done_pipe_write_req(0 downto 0),
      Block2_done_pipe_write_ack => Block2_done_pipe_write_ack(0 downto 0),
      Block2_done_pipe_write_data => Block2_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeC_tag_in,
      tag_out => convTransposeC_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeC_tag_in <= (others => '0');
  convTransposeC_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeC_start_req, start_ack => convTransposeC_start_ack,  fin_req => convTransposeC_fin_req,  fin_ack => convTransposeC_fin_ack);
  -- module convTransposeD
  convTransposeD_instance:convTransposeD-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeD_start_req,
      start_ack => convTransposeD_start_ack,
      fin_req => convTransposeD_fin_req,
      fin_ack => convTransposeD_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(18 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(0 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(0 downto 0),
      memory_space_3_sr_ack => memory_space_3_sr_ack(0 downto 0),
      memory_space_3_sr_addr => memory_space_3_sr_addr(13 downto 0),
      memory_space_3_sr_data => memory_space_3_sr_data(63 downto 0),
      memory_space_3_sr_tag => memory_space_3_sr_tag(18 downto 0),
      memory_space_3_sc_req => memory_space_3_sc_req(0 downto 0),
      memory_space_3_sc_ack => memory_space_3_sc_ack(0 downto 0),
      memory_space_3_sc_tag => memory_space_3_sc_tag(0 downto 0),
      Block1_start_pipe_read_req => Block1_start_pipe_read_req(0 downto 0),
      Block1_start_pipe_read_ack => Block1_start_pipe_read_ack(0 downto 0),
      Block1_start_pipe_read_data => Block1_start_pipe_read_data(15 downto 0),
      Block3_done_pipe_write_req => Block3_done_pipe_write_req(0 downto 0),
      Block3_done_pipe_write_ack => Block3_done_pipe_write_ack(0 downto 0),
      Block3_done_pipe_write_data => Block3_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeD_tag_in,
      tag_out => convTransposeD_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeD_tag_in <= (others => '0');
  convTransposeD_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeD_start_req, start_ack => convTransposeD_start_ack,  fin_req => convTransposeD_fin_req,  fin_ack => convTransposeD_fin_ack);
  -- module timer
  timer_out_args <= timer_c ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      c => timer_c,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(0 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(0 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  Block0_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_done_pipe_read_req,
      read_ack => Block0_done_pipe_read_ack,
      read_data => Block0_done_pipe_read_data,
      write_req => Block0_done_pipe_write_req,
      write_ack => Block0_done_pipe_write_ack,
      write_data => Block0_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block0_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_start_pipe_read_req,
      read_ack => Block0_start_pipe_read_ack,
      read_data => Block0_start_pipe_read_data,
      write_req => Block0_start_pipe_write_req,
      write_ack => Block0_start_pipe_write_ack,
      write_data => Block0_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_done_pipe_read_req,
      read_ack => Block1_done_pipe_read_ack,
      read_data => Block1_done_pipe_read_data,
      write_req => Block1_done_pipe_write_req,
      write_ack => Block1_done_pipe_write_ack,
      write_data => Block1_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_start",
      num_reads => 3,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_start_pipe_read_req,
      read_ack => Block1_start_pipe_read_ack,
      read_data => Block1_start_pipe_read_data,
      write_req => Block1_start_pipe_write_req,
      write_ack => Block1_start_pipe_write_ack,
      write_data => Block1_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_done_pipe_read_req,
      read_ack => Block2_done_pipe_read_ack,
      read_data => Block2_done_pipe_read_data,
      write_req => Block2_done_pipe_write_req,
      write_ack => Block2_done_pipe_write_ack,
      write_data => Block2_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_start_pipe_read_req,
      read_ack => Block2_start_pipe_read_ack,
      read_data => Block2_start_pipe_read_data,
      write_req => Block2_start_pipe_write_req,
      write_ack => Block2_start_pipe_write_ack,
      write_data => Block2_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_done_pipe_read_req,
      read_ack => Block3_done_pipe_read_ack,
      read_data => Block3_done_pipe_read_data,
      write_req => Block3_done_pipe_write_req,
      write_ack => Block3_done_pipe_write_ack,
      write_data => Block3_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_start_pipe_read_req,
      read_ack => Block3_start_pipe_read_ack,
      read_data => Block3_start_pipe_read_data,
      write_req => Block3_start_pipe_write_req,
      write_ack => Block3_start_pipe_write_ack,
      write_data => Block3_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_input_pipe_pipe_read_req,
      read_ack => ConvTranspose_input_pipe_pipe_read_ack,
      read_data => ConvTranspose_input_pipe_pipe_read_data,
      write_req => ConvTranspose_input_pipe_pipe_write_req,
      write_ack => ConvTranspose_input_pipe_pipe_write_ack,
      write_data => ConvTranspose_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_output_pipe_pipe_read_req,
      read_ack => ConvTranspose_output_pipe_pipe_read_ack,
      read_data => ConvTranspose_output_pipe_pipe_read_data,
      write_req => ConvTranspose_output_pipe_pipe_write_req,
      write_ack => ConvTranspose_output_pipe_pipe_write_ack,
      write_data => ConvTranspose_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  elapsed_time_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe elapsed_time_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => elapsed_time_pipe_pipe_read_req,
      read_ack => elapsed_time_pipe_pipe_read_ack,
      read_data => elapsed_time_pipe_pipe_read_data,
      write_req => elapsed_time_pipe_pipe_write_req,
      write_ack => elapsed_time_pipe_pipe_write_ack,
      write_data => elapsed_time_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  dummyROM_memory_space_0: dummy_read_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      addr_width => 1,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 4,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_2: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_stores => 1,
      addr_width => 11,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_3: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_3",
      num_loads => 1,
      num_stores => 5,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_3_lr_addr,
      lr_req_in => memory_space_3_lr_req,
      lr_ack_out => memory_space_3_lr_ack,
      lr_tag_in => memory_space_3_lr_tag,
      lc_req_in => memory_space_3_lc_req,
      lc_ack_out => memory_space_3_lc_ack,
      lc_data_out => memory_space_3_lc_data,
      lc_tag_out => memory_space_3_lc_tag,
      sr_addr_in => memory_space_3_sr_addr,
      sr_data_in => memory_space_3_sr_data,
      sr_req_in => memory_space_3_sr_req,
      sr_ack_out => memory_space_3_sr_ack,
      sr_tag_in => memory_space_3_sr_tag,
      sc_req_in=> memory_space_3_sc_req,
      sc_ack_out => memory_space_3_sc_ack,
      sc_tag_out => memory_space_3_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
