-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity fill_T is -- 
  generic (tag_length : integer); 
  port ( -- 
    addr : in  std_logic_vector(63 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(255 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(2 downto 0);
    maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity fill_T;
architecture fill_T_arch of fill_T is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal addr_buffer :  std_logic_vector(63 downto 0);
  signal addr_update_enable: Boolean;
  -- output port buffer signals
  signal fill_T_CP_0_start: Boolean;
  signal fill_T_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_maxpool_input_pipe_37_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_33_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_33_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_33_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_33_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_37_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_37_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_37_inst_ack_1 : boolean;
  signal CONCAT_u8_u16_38_inst_req_0 : boolean;
  signal CONCAT_u8_u16_38_inst_ack_0 : boolean;
  signal CONCAT_u8_u16_38_inst_req_1 : boolean;
  signal CONCAT_u8_u16_38_inst_ack_1 : boolean;
  signal CONCAT_u240_u256_45_inst_req_0 : boolean;
  signal CONCAT_u240_u256_45_inst_ack_0 : boolean;
  signal CONCAT_u240_u256_45_inst_req_1 : boolean;
  signal CONCAT_u240_u256_45_inst_ack_1 : boolean;
  signal addr_of_61_final_reg_ack_0 : boolean;
  signal addr_of_61_final_reg_req_1 : boolean;
  signal addr_of_61_final_reg_ack_1 : boolean;
  signal if_stmt_47_branch_req_0 : boolean;
  signal if_stmt_47_branch_ack_1 : boolean;
  signal if_stmt_47_branch_ack_0 : boolean;
  signal phi_stmt_15_req_1 : boolean;
  signal phi_stmt_21_req_1 : boolean;
  signal nmycount_31_17_buf_req_0 : boolean;
  signal nmycount_31_17_buf_ack_0 : boolean;
  signal nmycount_31_17_buf_req_1 : boolean;
  signal nmycount_31_17_buf_ack_1 : boolean;
  signal phi_stmt_15_req_0 : boolean;
  signal ninput_word_46_23_buf_req_0 : boolean;
  signal ninput_word_46_23_buf_ack_0 : boolean;
  signal ninput_word_46_23_buf_req_1 : boolean;
  signal ninput_word_46_23_buf_ack_1 : boolean;
  signal phi_stmt_21_req_0 : boolean;
  signal phi_stmt_15_ack_0 : boolean;
  signal phi_stmt_21_ack_0 : boolean;
  signal array_obj_ref_60_index_offset_req_0 : boolean;
  signal array_obj_ref_60_index_offset_ack_0 : boolean;
  signal array_obj_ref_60_index_offset_req_1 : boolean;
  signal array_obj_ref_60_index_offset_ack_1 : boolean;
  signal addr_of_61_final_reg_req_0 : boolean;
  signal ptr_deref_64_store_0_req_0 : boolean;
  signal ptr_deref_64_store_0_ack_0 : boolean;
  signal ptr_deref_64_store_0_req_1 : boolean;
  signal ptr_deref_64_store_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "fill_T_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 64) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(63 downto 0) <= addr;
  addr_buffer <= in_buffer_data_out(63 downto 0);
  in_buffer_data_in(tag_length + 63 downto 64) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 63 downto 64);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  fill_T_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "fill_T_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= fill_T_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= fill_T_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= fill_T_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  fill_T_CP_0: Block -- control-path 
    signal fill_T_CP_0_elements: BooleanArray(33 downto 0);
    -- 
  begin -- 
    fill_T_CP_0_elements(0) <= fill_T_CP_0_start;
    fill_T_CP_0_symbol <= fill_T_CP_0_elements(33);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	12 
    -- CP-element group 0:  members (5) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_13/$entry
      -- CP-element group 0: 	 branch_block_stmt_13/branch_block_stmt_13__entry__
      -- CP-element group 0: 	 branch_block_stmt_13/merge_stmt_14__entry__
      -- CP-element group 0: 	 branch_block_stmt_13/merge_stmt_14_dead_link/$entry
      -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	26 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	9 
    -- CP-element group 1: 	7 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (12) 
      -- CP-element group 1: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46__entry__
      -- CP-element group 1: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/$entry
      -- CP-element group 1: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_33_sample_start_
      -- CP-element group 1: 	 branch_block_stmt_13/merge_stmt_14__exit__
      -- CP-element group 1: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u8_u16_38_update_start_
      -- CP-element group 1: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_33_Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_33_Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u8_u16_38_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u8_u16_38_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u240_u256_45_update_start_
      -- CP-element group 1: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u240_u256_45_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u240_u256_45_Update/cr
      -- 
    rr_24_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_24_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(1), ack => RPIPE_maxpool_input_pipe_33_inst_req_0); -- 
    cr_57_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_57_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(1), ack => CONCAT_u8_u16_38_inst_req_1); -- 
    cr_71_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_71_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(1), ack => CONCAT_u240_u256_45_inst_req_1); -- 
    fill_T_CP_0_elements(1) <= fill_T_CP_0_elements(26);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_33_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_33_update_start_
      -- CP-element group 2: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_33_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_33_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_33_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_33_Update/cr
      -- 
    ra_25_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_33_inst_ack_0, ack => fill_T_CP_0_elements(2)); -- 
    cr_29_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_29_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(2), ack => RPIPE_maxpool_input_pipe_33_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_37_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_37_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_37_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_33_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_33_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_33_Update/ca
      -- 
    ca_30_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_33_inst_ack_1, ack => fill_T_CP_0_elements(3)); -- 
    rr_42_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_42_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(3), ack => RPIPE_maxpool_input_pipe_37_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_37_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_37_update_start_
      -- CP-element group 4: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_37_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_37_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_37_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_37_Update/cr
      -- 
    ra_43_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_37_inst_ack_0, ack => fill_T_CP_0_elements(4)); -- 
    cr_47_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_47_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(4), ack => RPIPE_maxpool_input_pipe_37_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u8_u16_38_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_37_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_37_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_37_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u8_u16_38_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u8_u16_38_Sample/rr
      -- 
    ca_48_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_37_inst_ack_1, ack => fill_T_CP_0_elements(5)); -- 
    rr_52_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_52_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(5), ack => CONCAT_u8_u16_38_inst_req_0); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u8_u16_38_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u8_u16_38_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u8_u16_38_Sample/ra
      -- 
    ra_53_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u8_u16_38_inst_ack_0, ack => fill_T_CP_0_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	1 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u8_u16_38_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u8_u16_38_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u8_u16_38_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u240_u256_45_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u240_u256_45_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u240_u256_45_Sample/rr
      -- 
    ca_58_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u8_u16_38_inst_ack_1, ack => fill_T_CP_0_elements(7)); -- 
    rr_66_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_66_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(7), ack => CONCAT_u240_u256_45_inst_req_0); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u240_u256_45_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u240_u256_45_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u240_u256_45_Sample/ra
      -- 
    ra_67_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u240_u256_45_inst_ack_0, ack => fill_T_CP_0_elements(8)); -- 
    -- CP-element group 9:  branch  transition  place  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	1 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (27) 
      -- CP-element group 9: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46__exit__
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47__entry__
      -- CP-element group 9: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/$exit
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47_eval_test/ULT_u4_u1_50/SplitProtocol/$entry
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47_eval_test/ULT_u4_u1_50/SplitProtocol/$exit
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47_eval_test/ULT_u4_u1_50/SplitProtocol/Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47_eval_test/ULT_u4_u1_50/SplitProtocol/Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u240_u256_45_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u240_u256_45_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u240_u256_45_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47_dead_link/$entry
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47_eval_test/$entry
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47_eval_test/$exit
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47_eval_test/ULT_u4_u1_50/$entry
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47_eval_test/ULT_u4_u1_50/$exit
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47_eval_test/ULT_u4_u1_50/ULT_u4_u1_50_inputs/$entry
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47_eval_test/ULT_u4_u1_50/ULT_u4_u1_50_inputs/$exit
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47_eval_test/ULT_u4_u1_50/SplitProtocol/Sample/rr
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47_eval_test/ULT_u4_u1_50/SplitProtocol/Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47_eval_test/ULT_u4_u1_50/SplitProtocol/Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47_eval_test/ULT_u4_u1_50/SplitProtocol/Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47_eval_test/ULT_u4_u1_50/SplitProtocol/Update/cr
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47_eval_test/ULT_u4_u1_50/SplitProtocol/Update/ca
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47_eval_test/branch_req
      -- CP-element group 9: 	 branch_block_stmt_13/ULT_u4_u1_50_place
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47_if_link/$entry
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47_else_link/$entry
      -- 
    ca_72_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u240_u256_45_inst_ack_1, ack => fill_T_CP_0_elements(9)); -- 
    branch_req_99_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_99_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(9), ack => if_stmt_47_branch_req_0); -- 
    -- CP-element group 10:  fork  transition  place  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	19 
    -- CP-element group 10: 	20 
    -- CP-element group 10: 	17 
    -- CP-element group 10: 	16 
    -- CP-element group 10:  members (18) 
      -- CP-element group 10: 	 branch_block_stmt_13/if_stmt_47_if_link/$exit
      -- CP-element group 10: 	 branch_block_stmt_13/if_stmt_47_if_link/if_choice_transition
      -- CP-element group 10: 	 branch_block_stmt_13/loopback
      -- CP-element group 10: 	 branch_block_stmt_13/loopback_PhiReq/$entry
      -- CP-element group 10: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_15/$entry
      -- CP-element group 10: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_15/phi_stmt_15_sources/$entry
      -- CP-element group 10: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_15/phi_stmt_15_sources/Interlock/$entry
      -- CP-element group 10: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_15/phi_stmt_15_sources/Interlock/Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_15/phi_stmt_15_sources/Interlock/Sample/req
      -- CP-element group 10: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_15/phi_stmt_15_sources/Interlock/Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_15/phi_stmt_15_sources/Interlock/Update/req
      -- CP-element group 10: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_21/$entry
      -- CP-element group 10: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_21/phi_stmt_21_sources/$entry
      -- CP-element group 10: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_21/phi_stmt_21_sources/Interlock/$entry
      -- CP-element group 10: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_21/phi_stmt_21_sources/Interlock/Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_21/phi_stmt_21_sources/Interlock/Sample/req
      -- CP-element group 10: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_21/phi_stmt_21_sources/Interlock/Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_21/phi_stmt_21_sources/Interlock/Update/req
      -- 
    if_choice_transition_104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_47_branch_ack_1, ack => fill_T_CP_0_elements(10)); -- 
    req_148_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_148_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(10), ack => nmycount_31_17_buf_req_0); -- 
    req_153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(10), ack => nmycount_31_17_buf_req_1); -- 
    req_168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(10), ack => ninput_word_46_23_buf_req_0); -- 
    req_173_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_173_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(10), ack => ninput_word_46_23_buf_req_1); -- 
    -- CP-element group 11:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	27 
    -- CP-element group 11: 	28 
    -- CP-element group 11: 	30 
    -- CP-element group 11: 	32 
    -- CP-element group 11:  members (30) 
      -- CP-element group 11: 	 branch_block_stmt_13/branch_block_stmt_13__exit__
      -- CP-element group 11: 	 branch_block_stmt_13/if_stmt_47__exit__
      -- CP-element group 11: 	 branch_block_stmt_13/$exit
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/addr_of_61_complete/$entry
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/addr_of_61_complete/req
      -- CP-element group 11: 	 branch_block_stmt_13/if_stmt_47_else_link/$exit
      -- CP-element group 11: 	 branch_block_stmt_13/if_stmt_47_else_link/else_choice_transition
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/$entry
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/addr_of_61_update_start_
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_index_resized_1
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_index_scaled_1
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_index_computed_1
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_index_resize_1/$entry
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_index_resize_1/$exit
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_index_resize_1/index_resize_req
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_index_resize_1/index_resize_ack
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_index_scale_1/$entry
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_index_scale_1/$exit
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_index_scale_1/scale_rename_req
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_index_scale_1/scale_rename_ack
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_final_index_sum_regn_update_start
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_final_index_sum_regn_Sample/$entry
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_final_index_sum_regn_Sample/req
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_final_index_sum_regn_Update/$entry
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_final_index_sum_regn_Update/req
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_update_start_
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_Update/$entry
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_Update/word_access_complete/$entry
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_Update/word_access_complete/word_0/$entry
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_Update/word_access_complete/word_0/cr
      -- 
    else_choice_transition_108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_47_branch_ack_0, ack => fill_T_CP_0_elements(11)); -- 
    req_229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(11), ack => addr_of_61_final_reg_req_1); -- 
    req_209_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_209_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(11), ack => array_obj_ref_60_index_offset_req_0); -- 
    req_214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(11), ack => array_obj_ref_60_index_offset_req_1); -- 
    cr_279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(11), ack => ptr_deref_64_store_0_req_1); -- 
    -- CP-element group 12:  fork  transition  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	14 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (5) 
      -- CP-element group 12: 	 branch_block_stmt_13/merge_stmt_14__entry___PhiReq/$entry
      -- CP-element group 12: 	 branch_block_stmt_13/merge_stmt_14__entry___PhiReq/phi_stmt_15/$entry
      -- CP-element group 12: 	 branch_block_stmt_13/merge_stmt_14__entry___PhiReq/phi_stmt_15/phi_stmt_15_sources/$entry
      -- CP-element group 12: 	 branch_block_stmt_13/merge_stmt_14__entry___PhiReq/phi_stmt_21/$entry
      -- CP-element group 12: 	 branch_block_stmt_13/merge_stmt_14__entry___PhiReq/phi_stmt_21/phi_stmt_21_sources/$entry
      -- 
    fill_T_CP_0_elements(12) <= fill_T_CP_0_elements(0);
    -- CP-element group 13:  transition  output  delay-element  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	15 
    -- CP-element group 13:  members (4) 
      -- CP-element group 13: 	 branch_block_stmt_13/merge_stmt_14__entry___PhiReq/phi_stmt_15/$exit
      -- CP-element group 13: 	 branch_block_stmt_13/merge_stmt_14__entry___PhiReq/phi_stmt_15/phi_stmt_15_sources/$exit
      -- CP-element group 13: 	 branch_block_stmt_13/merge_stmt_14__entry___PhiReq/phi_stmt_15/phi_stmt_15_sources/type_cast_20_konst_delay_trans
      -- CP-element group 13: 	 branch_block_stmt_13/merge_stmt_14__entry___PhiReq/phi_stmt_15/phi_stmt_15_req
      -- 
    phi_stmt_15_req_124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_15_req_124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(13), ack => phi_stmt_15_req_1); -- 
    -- Element group fill_T_CP_0_elements(13) is a control-delay.
    cp_element_13_delay: control_delay_element  generic map(name => " 13_delay", delay_value => 1)  port map(req => fill_T_CP_0_elements(12), ack => fill_T_CP_0_elements(13), clk => clk, reset =>reset);
    -- CP-element group 14:  transition  output  delay-element  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	12 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (4) 
      -- CP-element group 14: 	 branch_block_stmt_13/merge_stmt_14__entry___PhiReq/phi_stmt_21/$exit
      -- CP-element group 14: 	 branch_block_stmt_13/merge_stmt_14__entry___PhiReq/phi_stmt_21/phi_stmt_21_sources/$exit
      -- CP-element group 14: 	 branch_block_stmt_13/merge_stmt_14__entry___PhiReq/phi_stmt_21/phi_stmt_21_sources/type_cast_25_konst_delay_trans
      -- CP-element group 14: 	 branch_block_stmt_13/merge_stmt_14__entry___PhiReq/phi_stmt_21/phi_stmt_21_req
      -- 
    phi_stmt_21_req_132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_21_req_132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(14), ack => phi_stmt_21_req_1); -- 
    -- Element group fill_T_CP_0_elements(14) is a control-delay.
    cp_element_14_delay: control_delay_element  generic map(name => " 14_delay", delay_value => 1)  port map(req => fill_T_CP_0_elements(12), ack => fill_T_CP_0_elements(14), clk => clk, reset =>reset);
    -- CP-element group 15:  join  transition  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: 	13 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	23 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_13/merge_stmt_14__entry___PhiReq/$exit
      -- 
    fill_T_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "fill_T_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= fill_T_CP_0_elements(14) & fill_T_CP_0_elements(13);
      gj_fill_T_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => fill_T_CP_0_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	10 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	18 
    -- CP-element group 16:  members (2) 
      -- CP-element group 16: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_15/phi_stmt_15_sources/Interlock/Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_15/phi_stmt_15_sources/Interlock/Sample/ack
      -- 
    ack_149_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_31_17_buf_ack_0, ack => fill_T_CP_0_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	10 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_15/phi_stmt_15_sources/Interlock/Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_15/phi_stmt_15_sources/Interlock/Update/ack
      -- 
    ack_154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_31_17_buf_ack_1, ack => fill_T_CP_0_elements(17)); -- 
    -- CP-element group 18:  join  transition  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: 	16 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	22 
    -- CP-element group 18:  members (4) 
      -- CP-element group 18: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_15/$exit
      -- CP-element group 18: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_15/phi_stmt_15_sources/$exit
      -- CP-element group 18: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_15/phi_stmt_15_sources/Interlock/$exit
      -- CP-element group 18: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_15/phi_stmt_15_req
      -- 
    phi_stmt_15_req_155_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_15_req_155_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(18), ack => phi_stmt_15_req_0); -- 
    fill_T_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "fill_T_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= fill_T_CP_0_elements(17) & fill_T_CP_0_elements(16);
      gj_fill_T_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => fill_T_CP_0_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	10 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	21 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_21/phi_stmt_21_sources/Interlock/Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_21/phi_stmt_21_sources/Interlock/Sample/ack
      -- 
    ack_169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ninput_word_46_23_buf_ack_0, ack => fill_T_CP_0_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	10 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_21/phi_stmt_21_sources/Interlock/Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_21/phi_stmt_21_sources/Interlock/Update/ack
      -- 
    ack_174_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ninput_word_46_23_buf_ack_1, ack => fill_T_CP_0_elements(20)); -- 
    -- CP-element group 21:  join  transition  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	19 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (4) 
      -- CP-element group 21: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_21/$exit
      -- CP-element group 21: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_21/phi_stmt_21_sources/$exit
      -- CP-element group 21: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_21/phi_stmt_21_sources/Interlock/$exit
      -- CP-element group 21: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_21/phi_stmt_21_req
      -- 
    phi_stmt_21_req_175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_21_req_175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(21), ack => phi_stmt_21_req_0); -- 
    fill_T_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "fill_T_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= fill_T_CP_0_elements(19) & fill_T_CP_0_elements(20);
      gj_fill_T_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => fill_T_CP_0_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  transition  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: 	18 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_13/loopback_PhiReq/$exit
      -- 
    fill_T_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "fill_T_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= fill_T_CP_0_elements(21) & fill_T_CP_0_elements(18);
      gj_fill_T_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => fill_T_CP_0_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  merge  fork  transition  place  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: 	15 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	25 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_13/merge_stmt_14_PhiReqMerge
      -- CP-element group 23: 	 branch_block_stmt_13/merge_stmt_14_PhiAck/$entry
      -- 
    fill_T_CP_0_elements(23) <= OrReduce(fill_T_CP_0_elements(22) & fill_T_CP_0_elements(15));
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_13/merge_stmt_14_PhiAck/phi_stmt_15_ack
      -- 
    phi_stmt_15_ack_180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_15_ack_0, ack => fill_T_CP_0_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	23 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_13/merge_stmt_14_PhiAck/phi_stmt_21_ack
      -- 
    phi_stmt_21_ack_181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_21_ack_0, ack => fill_T_CP_0_elements(25)); -- 
    -- CP-element group 26:  join  transition  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	1 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_13/merge_stmt_14_PhiAck/$exit
      -- 
    fill_T_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "fill_T_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= fill_T_CP_0_elements(25) & fill_T_CP_0_elements(24);
      gj_fill_T_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => fill_T_CP_0_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	11 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	33 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_final_index_sum_regn_sample_complete
      -- CP-element group 27: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_final_index_sum_regn_Sample/$exit
      -- CP-element group 27: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_final_index_sum_regn_Sample/ack
      -- 
    ack_210_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_60_index_offset_ack_0, ack => fill_T_CP_0_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	11 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (11) 
      -- CP-element group 28: 	 assign_stmt_62_to_assign_stmt_66/addr_of_61_sample_start_
      -- CP-element group 28: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_root_address_calculated
      -- CP-element group 28: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_offset_calculated
      -- CP-element group 28: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_final_index_sum_regn_Update/$exit
      -- CP-element group 28: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_final_index_sum_regn_Update/ack
      -- CP-element group 28: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_base_plus_offset/$entry
      -- CP-element group 28: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_base_plus_offset/$exit
      -- CP-element group 28: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_base_plus_offset/sum_rename_req
      -- CP-element group 28: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_base_plus_offset/sum_rename_ack
      -- CP-element group 28: 	 assign_stmt_62_to_assign_stmt_66/addr_of_61_request/$entry
      -- CP-element group 28: 	 assign_stmt_62_to_assign_stmt_66/addr_of_61_request/req
      -- 
    ack_215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_60_index_offset_ack_1, ack => fill_T_CP_0_elements(28)); -- 
    req_224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(28), ack => addr_of_61_final_reg_req_0); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 assign_stmt_62_to_assign_stmt_66/addr_of_61_request/ack
      -- CP-element group 29: 	 assign_stmt_62_to_assign_stmt_66/addr_of_61_sample_completed_
      -- CP-element group 29: 	 assign_stmt_62_to_assign_stmt_66/addr_of_61_request/$exit
      -- 
    ack_225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_61_final_reg_ack_0, ack => fill_T_CP_0_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	11 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (28) 
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/addr_of_61_complete/$exit
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/addr_of_61_complete/ack
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/addr_of_61_update_completed_
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_sample_start_
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_base_address_calculated
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_word_address_calculated
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_root_address_calculated
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_base_address_resized
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_base_addr_resize/$entry
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_base_addr_resize/$exit
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_base_addr_resize/base_resize_req
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_base_addr_resize/base_resize_ack
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_base_plus_offset/$entry
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_base_plus_offset/$exit
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_base_plus_offset/sum_rename_req
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_base_plus_offset/sum_rename_ack
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_word_addrgen/$entry
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_word_addrgen/$exit
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_word_addrgen/root_register_req
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_word_addrgen/root_register_ack
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_Sample/$entry
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_Sample/ptr_deref_64_Split/$entry
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_Sample/ptr_deref_64_Split/$exit
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_Sample/ptr_deref_64_Split/split_req
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_Sample/ptr_deref_64_Split/split_ack
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_Sample/word_access_start/$entry
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_Sample/word_access_start/word_0/$entry
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_Sample/word_access_start/word_0/rr
      -- 
    ack_230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_61_final_reg_ack_1, ack => fill_T_CP_0_elements(30)); -- 
    rr_268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(30), ack => ptr_deref_64_store_0_req_0); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (5) 
      -- CP-element group 31: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_sample_completed_
      -- CP-element group 31: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_Sample/$exit
      -- CP-element group 31: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_Sample/word_access_start/$exit
      -- CP-element group 31: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_Sample/word_access_start/word_0/$exit
      -- CP-element group 31: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_Sample/word_access_start/word_0/ra
      -- 
    ra_269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_64_store_0_ack_0, ack => fill_T_CP_0_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	11 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (5) 
      -- CP-element group 32: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_update_completed_
      -- CP-element group 32: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_Update/$exit
      -- CP-element group 32: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_Update/word_access_complete/$exit
      -- CP-element group 32: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_Update/word_access_complete/word_0/$exit
      -- CP-element group 32: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_Update/word_access_complete/word_0/ca
      -- 
    ca_280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_64_store_0_ack_1, ack => fill_T_CP_0_elements(32)); -- 
    -- CP-element group 33:  join  transition  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	27 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (2) 
      -- CP-element group 33: 	 $exit
      -- CP-element group 33: 	 assign_stmt_62_to_assign_stmt_66/$exit
      -- 
    fill_T_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "fill_T_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= fill_T_CP_0_elements(27) & fill_T_CP_0_elements(32);
      gj_fill_T_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => fill_T_CP_0_elements(33), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal RPIPE_maxpool_input_pipe_37_wire : std_logic_vector(7 downto 0);
    signal R_addr_59_resized : std_logic_vector(13 downto 0);
    signal R_addr_59_scaled : std_logic_vector(13 downto 0);
    signal ULT_u4_u1_50_wire : std_logic_vector(0 downto 0);
    signal array_obj_ref_60_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_60_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_60_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_60_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_60_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_60_root_address : std_logic_vector(13 downto 0);
    signal input_word_21 : std_logic_vector(255 downto 0);
    signal konst_29_wire_constant : std_logic_vector(3 downto 0);
    signal konst_49_wire_constant : std_logic_vector(3 downto 0);
    signal mycount_15 : std_logic_vector(3 downto 0);
    signal ninput_word_46 : std_logic_vector(255 downto 0);
    signal ninput_word_46_23_buffered : std_logic_vector(255 downto 0);
    signal nmycount_31 : std_logic_vector(3 downto 0);
    signal nmycount_31_17_buffered : std_logic_vector(3 downto 0);
    signal ptr_62 : std_logic_vector(31 downto 0);
    signal ptr_deref_64_data_0 : std_logic_vector(255 downto 0);
    signal ptr_deref_64_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_64_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_64_wire : std_logic_vector(255 downto 0);
    signal ptr_deref_64_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_64_word_offset_0 : std_logic_vector(13 downto 0);
    signal slice_43_wire : std_logic_vector(239 downto 0);
    signal type_cast_20_wire_constant : std_logic_vector(3 downto 0);
    signal type_cast_25_wire_constant : std_logic_vector(255 downto 0);
    signal val1_34 : std_logic_vector(7 downto 0);
    signal val_39 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_60_constant_part_of_offset <= "00000000000000";
    array_obj_ref_60_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_60_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_60_resized_base_address <= "00000000000000";
    konst_29_wire_constant <= "0001";
    konst_49_wire_constant <= "1111";
    ptr_deref_64_word_offset_0 <= "00000000000000";
    type_cast_20_wire_constant <= "0000";
    type_cast_25_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_15: Block -- phi operator 
      signal idata: std_logic_vector(7 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nmycount_31_17_buffered & type_cast_20_wire_constant;
      req <= phi_stmt_15_req_0 & phi_stmt_15_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_15",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 4) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_15_ack_0,
          idata => idata,
          odata => mycount_15,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_15
    phi_stmt_21: Block -- phi operator 
      signal idata: std_logic_vector(511 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= ninput_word_46_23_buffered & type_cast_25_wire_constant;
      req <= phi_stmt_21_req_0 & phi_stmt_21_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_21",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 256) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_21_ack_0,
          idata => idata,
          odata => input_word_21,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_21
    -- flow-through slice operator slice_43_inst
    slice_43_wire <= input_word_21(239 downto 0);
    addr_of_61_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_61_final_reg_req_0;
      addr_of_61_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_61_final_reg_req_1;
      addr_of_61_final_reg_ack_1<= rack(0);
      addr_of_61_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_61_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_60_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ptr_62,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    ninput_word_46_23_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= ninput_word_46_23_buf_req_0;
      ninput_word_46_23_buf_ack_0<= wack(0);
      rreq(0) <= ninput_word_46_23_buf_req_1;
      ninput_word_46_23_buf_ack_1<= rack(0);
      ninput_word_46_23_buf : InterlockBuffer generic map ( -- 
        name => "ninput_word_46_23_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 256,
        out_data_width => 256,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ninput_word_46,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ninput_word_46_23_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nmycount_31_17_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nmycount_31_17_buf_req_0;
      nmycount_31_17_buf_ack_0<= wack(0);
      rreq(0) <= nmycount_31_17_buf_req_1;
      nmycount_31_17_buf_ack_1<= rack(0);
      nmycount_31_17_buf : InterlockBuffer generic map ( -- 
        name => "nmycount_31_17_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 4,
        out_data_width => 4,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nmycount_31,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nmycount_31_17_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_60_index_1_rename
    process(R_addr_59_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr_59_resized;
      ov(13 downto 0) := iv;
      R_addr_59_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_60_index_1_resize
    process(addr_buffer) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr_buffer;
      ov := iv(13 downto 0);
      R_addr_59_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_60_root_address_inst
    process(array_obj_ref_60_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_60_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_60_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_64_addr_0
    process(ptr_deref_64_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_64_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_64_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_64_base_resize
    process(ptr_62) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_62;
      ov := iv(13 downto 0);
      ptr_deref_64_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_64_gather_scatter
    process(ninput_word_46) --
      variable iv : std_logic_vector(255 downto 0);
      variable ov : std_logic_vector(255 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ninput_word_46;
      ov(255 downto 0) := iv;
      ptr_deref_64_data_0 <= ov(255 downto 0);
      --
    end process;
    -- equivalence ptr_deref_64_root_address_inst
    process(ptr_deref_64_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_64_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_64_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_47_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u4_u1_50_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_47_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_47_branch_req_0,
          ack0 => if_stmt_47_branch_ack_0,
          ack1 => if_stmt_47_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u4_u4_30_inst
    process(mycount_15) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mycount_15, konst_29_wire_constant, tmp_var);
      nmycount_31 <= tmp_var; --
    end process;
    -- shared split operator group (1) : CONCAT_u240_u256_45_inst 
    ApConcat_group_1: Block -- 
      signal data_in: std_logic_vector(255 downto 0);
      signal data_out: std_logic_vector(255 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= slice_43_wire & val_39;
      ninput_word_46 <= data_out(255 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u240_u256_45_inst_req_0;
      CONCAT_u240_u256_45_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u240_u256_45_inst_req_1;
      CONCAT_u240_u256_45_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_1_gI: SplitGuardInterface generic map(name => "ApConcat_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 240,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 256,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : CONCAT_u8_u16_38_inst 
    ApConcat_group_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= val1_34 & RPIPE_maxpool_input_pipe_37_wire;
      val_39 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u8_u16_38_inst_req_0;
      CONCAT_u8_u16_38_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u8_u16_38_inst_req_1;
      CONCAT_u8_u16_38_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_2_gI: SplitGuardInterface generic map(name => "ApConcat_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_2",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- binary operator ULT_u4_u1_50_inst
    process(mycount_15) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(mycount_15, konst_49_wire_constant, tmp_var);
      ULT_u4_u1_50_wire <= tmp_var; --
    end process;
    -- shared split operator group (4) : array_obj_ref_60_index_offset 
    ApIntAdd_group_4: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_addr_59_scaled;
      array_obj_ref_60_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_60_index_offset_req_0;
      array_obj_ref_60_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_60_index_offset_req_1;
      array_obj_ref_60_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_4_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_4",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared store operator group (0) : ptr_deref_64_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(255 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_64_store_0_req_0;
      ptr_deref_64_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_64_store_0_req_1;
      ptr_deref_64_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_64_word_address_0;
      data_in <= ptr_deref_64_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 256,
        num_reqs => 1,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(255 downto 0),
          mtag => memory_space_1_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_maxpool_input_pipe_33_inst RPIPE_maxpool_input_pipe_37_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 1 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= RPIPE_maxpool_input_pipe_33_inst_req_0;
      reqL_unguarded(0) <= RPIPE_maxpool_input_pipe_37_inst_req_0;
      RPIPE_maxpool_input_pipe_33_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_maxpool_input_pipe_37_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= RPIPE_maxpool_input_pipe_33_inst_req_1;
      reqR_unguarded(0) <= RPIPE_maxpool_input_pipe_37_inst_req_1;
      RPIPE_maxpool_input_pipe_33_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_maxpool_input_pipe_37_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      val1_34 <= data_out(15 downto 8);
      RPIPE_maxpool_input_pipe_37_wire <= data_out(7 downto 0);
      maxpool_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "maxpool_input_pipe_read_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      maxpool_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "maxpool_input_pipe_read_0", data_width => 8,  num_reqs => 2,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => maxpool_input_pipe_pipe_read_req(0),
          oack => maxpool_input_pipe_pipe_read_ack(0),
          odata => maxpool_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- 
  end Block; -- data_path
  -- 
end fill_T_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity maxPool3D is -- 
  generic (tag_length : integer); 
  port ( -- 
    maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    fill_T_call_reqs : out  std_logic_vector(0 downto 0);
    fill_T_call_acks : in   std_logic_vector(0 downto 0);
    fill_T_call_data : out  std_logic_vector(63 downto 0);
    fill_T_call_tag  :  out  std_logic_vector(0 downto 0);
    fill_T_return_reqs : out  std_logic_vector(0 downto 0);
    fill_T_return_acks : in   std_logic_vector(0 downto 0);
    fill_T_return_tag :  in   std_logic_vector(0 downto 0);
    maxPool4_call_reqs : out  std_logic_vector(0 downto 0);
    maxPool4_call_acks : in   std_logic_vector(0 downto 0);
    maxPool4_call_data : out  std_logic_vector(159 downto 0);
    maxPool4_call_tag  :  out  std_logic_vector(0 downto 0);
    maxPool4_return_reqs : out  std_logic_vector(0 downto 0);
    maxPool4_return_acks : in   std_logic_vector(0 downto 0);
    maxPool4_return_data : in   std_logic_vector(7 downto 0);
    maxPool4_return_tag :  in   std_logic_vector(0 downto 0);
    sendB_call_reqs : out  std_logic_vector(0 downto 0);
    sendB_call_acks : in   std_logic_vector(0 downto 0);
    sendB_call_data : out  std_logic_vector(31 downto 0);
    sendB_call_tag  :  out  std_logic_vector(0 downto 0);
    sendB_return_reqs : out  std_logic_vector(0 downto 0);
    sendB_return_acks : in   std_logic_vector(0 downto 0);
    sendB_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity maxPool3D;
architecture maxPool3D_arch of maxPool3D is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal maxPool3D_CP_2619_start: Boolean;
  signal maxPool3D_CP_2619_symbol: Boolean;
  -- volatile/operator module components. 
  component fill_T is -- 
    generic (tag_length : integer); 
    port ( -- 
      addr : in  std_logic_vector(63 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(255 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(2 downto 0);
      maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component maxPool4 is -- 
    generic (tag_length : integer); 
    port ( -- 
      addr : in  std_logic_vector(31 downto 0);
      addr1 : in  std_logic_vector(31 downto 0);
      addr2 : in  std_logic_vector(31 downto 0);
      addr3 : in  std_logic_vector(31 downto 0);
      addr4 : in  std_logic_vector(31 downto 0);
      output : out  std_logic_vector(7 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(255 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component sendB is -- 
    generic (tag_length : integer); 
    port ( -- 
      size : in  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal type_cast_1346_inst_ack_1 : boolean;
  signal type_cast_1830_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1367_inst_ack_1 : boolean;
  signal type_cast_1346_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1392_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1367_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1354_inst_ack_0 : boolean;
  signal type_cast_1383_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1379_inst_req_0 : boolean;
  signal type_cast_1358_inst_ack_1 : boolean;
  signal type_cast_1358_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1404_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1379_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1329_inst_req_0 : boolean;
  signal call_stmt_1743_call_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1404_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1392_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1392_inst_req_0 : boolean;
  signal type_cast_1383_inst_ack_1 : boolean;
  signal type_cast_1333_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1329_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1417_inst_req_0 : boolean;
  signal type_cast_1396_inst_req_1 : boolean;
  signal type_cast_1656_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1354_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1392_inst_ack_1 : boolean;
  signal type_cast_1661_inst_req_1 : boolean;
  signal call_stmt_1743_call_ack_0 : boolean;
  signal type_cast_1396_inst_req_0 : boolean;
  signal call_stmt_1743_call_req_0 : boolean;
  signal call_stmt_1743_call_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1815_inst_ack_1 : boolean;
  signal W_colx_x1_1749_delayed_1_0_1759_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1329_inst_req_1 : boolean;
  signal type_cast_1396_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1354_inst_ack_1 : boolean;
  signal type_cast_1661_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1329_inst_ack_1 : boolean;
  signal W_colx_x1_1749_delayed_1_0_1759_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1404_inst_req_0 : boolean;
  signal type_cast_1371_inst_ack_1 : boolean;
  signal type_cast_1333_inst_req_1 : boolean;
  signal type_cast_1371_inst_req_1 : boolean;
  signal type_cast_1757_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1354_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1367_inst_ack_0 : boolean;
  signal type_cast_1346_inst_ack_0 : boolean;
  signal type_cast_1358_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1342_inst_ack_1 : boolean;
  signal type_cast_1358_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1342_inst_req_1 : boolean;
  signal type_cast_1757_inst_req_0 : boolean;
  signal type_cast_1830_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1367_inst_req_0 : boolean;
  signal type_cast_1559_inst_req_1 : boolean;
  signal type_cast_1346_inst_req_0 : boolean;
  signal phi_stmt_1553_ack_0 : boolean;
  signal type_cast_1371_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1342_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1379_inst_ack_1 : boolean;
  signal type_cast_1559_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1342_inst_req_0 : boolean;
  signal type_cast_1371_inst_req_0 : boolean;
  signal type_cast_1826_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1379_inst_req_1 : boolean;
  signal type_cast_1333_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1404_inst_ack_0 : boolean;
  signal type_cast_1559_inst_req_0 : boolean;
  signal type_cast_1383_inst_req_1 : boolean;
  signal type_cast_1383_inst_ack_0 : boolean;
  signal type_cast_1826_inst_ack_0 : boolean;
  signal type_cast_1333_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1815_inst_req_1 : boolean;
  signal type_cast_1559_inst_ack_1 : boolean;
  signal type_cast_1396_inst_ack_0 : boolean;
  signal phi_stmt_1553_req_1 : boolean;
  signal type_cast_1656_inst_req_1 : boolean;
  signal type_cast_1656_inst_ack_1 : boolean;
  signal type_cast_1408_inst_req_0 : boolean;
  signal type_cast_1408_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1815_inst_ack_0 : boolean;
  signal type_cast_1408_inst_req_1 : boolean;
  signal do_while_stmt_1646_branch_ack_1 : boolean;
  signal type_cast_1408_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1815_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1417_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1417_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1417_inst_ack_1 : boolean;
  signal type_cast_1674_inst_ack_1 : boolean;
  signal type_cast_1674_inst_req_1 : boolean;
  signal type_cast_1421_inst_req_0 : boolean;
  signal do_while_stmt_1646_branch_ack_0 : boolean;
  signal type_cast_1421_inst_ack_0 : boolean;
  signal type_cast_1421_inst_req_1 : boolean;
  signal type_cast_1421_inst_ack_1 : boolean;
  signal type_cast_1661_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1429_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1429_inst_ack_0 : boolean;
  signal type_cast_1661_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1429_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1429_inst_ack_1 : boolean;
  signal type_cast_1674_inst_ack_0 : boolean;
  signal type_cast_1674_inst_req_0 : boolean;
  signal W_rowx_x1_1770_delayed_2_0_1783_inst_ack_1 : boolean;
  signal type_cast_1433_inst_req_0 : boolean;
  signal W_rowx_x1_1770_delayed_2_0_1783_inst_req_1 : boolean;
  signal type_cast_1433_inst_ack_0 : boolean;
  signal type_cast_1433_inst_req_1 : boolean;
  signal type_cast_1433_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1442_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1442_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1442_inst_req_1 : boolean;
  signal W_rowx_x1_1770_delayed_2_0_1783_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1442_inst_ack_1 : boolean;
  signal type_cast_1670_inst_ack_1 : boolean;
  signal W_rowx_x1_1770_delayed_2_0_1783_inst_req_0 : boolean;
  signal call_stmt_1843_call_ack_1 : boolean;
  signal type_cast_1446_inst_req_0 : boolean;
  signal type_cast_1446_inst_ack_0 : boolean;
  signal call_stmt_1843_call_req_1 : boolean;
  signal type_cast_1446_inst_req_1 : boolean;
  signal type_cast_1446_inst_ack_1 : boolean;
  signal if_stmt_1809_branch_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1819_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1819_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1454_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1454_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1454_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1454_inst_ack_1 : boolean;
  signal type_cast_1670_inst_req_1 : boolean;
  signal type_cast_1458_inst_req_0 : boolean;
  signal type_cast_1458_inst_ack_0 : boolean;
  signal type_cast_1458_inst_req_1 : boolean;
  signal type_cast_1781_inst_ack_1 : boolean;
  signal type_cast_1458_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1819_inst_ack_0 : boolean;
  signal type_cast_1670_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1467_inst_req_0 : boolean;
  signal type_cast_1781_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1467_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1467_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1467_inst_ack_1 : boolean;
  signal type_cast_1670_inst_req_0 : boolean;
  signal phi_stmt_1553_req_0 : boolean;
  signal call_stmt_1843_call_ack_0 : boolean;
  signal type_cast_1471_inst_req_0 : boolean;
  signal type_cast_1471_inst_ack_0 : boolean;
  signal call_stmt_1843_call_req_0 : boolean;
  signal type_cast_1471_inst_req_1 : boolean;
  signal type_cast_1781_inst_ack_0 : boolean;
  signal type_cast_1471_inst_ack_1 : boolean;
  signal if_stmt_1809_branch_ack_1 : boolean;
  signal type_cast_1826_inst_ack_1 : boolean;
  signal type_cast_1826_inst_req_1 : boolean;
  signal type_cast_1666_inst_ack_1 : boolean;
  signal type_cast_1781_inst_req_0 : boolean;
  signal type_cast_1666_inst_req_1 : boolean;
  signal type_cast_1481_inst_req_0 : boolean;
  signal type_cast_1481_inst_ack_0 : boolean;
  signal type_cast_1656_inst_req_0 : boolean;
  signal type_cast_1481_inst_req_1 : boolean;
  signal type_cast_1481_inst_ack_1 : boolean;
  signal phi_stmt_1658_ack_0 : boolean;
  signal if_stmt_1499_branch_req_0 : boolean;
  signal type_cast_1757_inst_ack_1 : boolean;
  signal if_stmt_1499_branch_ack_1 : boolean;
  signal if_stmt_1499_branch_ack_0 : boolean;
  signal type_cast_1757_inst_req_1 : boolean;
  signal type_cast_1666_inst_ack_0 : boolean;
  signal type_cast_1536_inst_req_0 : boolean;
  signal type_cast_1536_inst_ack_0 : boolean;
  signal type_cast_1536_inst_req_1 : boolean;
  signal type_cast_1536_inst_ack_1 : boolean;
  signal phi_stmt_1658_req_1 : boolean;
  signal type_cast_1666_inst_req_0 : boolean;
  signal type_cast_1830_inst_ack_1 : boolean;
  signal call_stmt_1562_call_req_0 : boolean;
  signal W_colx_x1_1749_delayed_1_0_1759_inst_ack_1 : boolean;
  signal call_stmt_1562_call_ack_0 : boolean;
  signal type_cast_1830_inst_req_1 : boolean;
  signal call_stmt_1562_call_req_1 : boolean;
  signal W_colx_x1_1749_delayed_1_0_1759_inst_req_1 : boolean;
  signal call_stmt_1562_call_ack_1 : boolean;
  signal if_stmt_1809_branch_req_0 : boolean;
  signal phi_stmt_1658_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1819_inst_req_0 : boolean;
  signal if_stmt_1574_branch_req_0 : boolean;
  signal if_stmt_1574_branch_ack_1 : boolean;
  signal if_stmt_1574_branch_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1596_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1596_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1596_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1596_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1600_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1600_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1600_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1600_inst_ack_1 : boolean;
  signal type_cast_1607_inst_req_0 : boolean;
  signal type_cast_1607_inst_ack_0 : boolean;
  signal type_cast_1607_inst_req_1 : boolean;
  signal type_cast_1607_inst_ack_1 : boolean;
  signal type_cast_1611_inst_req_0 : boolean;
  signal type_cast_1611_inst_ack_0 : boolean;
  signal type_cast_1611_inst_req_1 : boolean;
  signal type_cast_1611_inst_ack_1 : boolean;
  signal type_cast_1615_inst_req_0 : boolean;
  signal type_cast_1615_inst_ack_0 : boolean;
  signal type_cast_1615_inst_req_1 : boolean;
  signal type_cast_1615_inst_ack_1 : boolean;
  signal do_while_stmt_1646_branch_req_0 : boolean;
  signal phi_stmt_1648_req_0 : boolean;
  signal phi_stmt_1648_req_1 : boolean;
  signal phi_stmt_1648_ack_0 : boolean;
  signal type_cast_1651_inst_req_0 : boolean;
  signal type_cast_1651_inst_ack_0 : boolean;
  signal type_cast_1651_inst_req_1 : boolean;
  signal type_cast_1651_inst_ack_1 : boolean;
  signal phi_stmt_1653_req_0 : boolean;
  signal phi_stmt_1653_req_1 : boolean;
  signal phi_stmt_1653_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "maxPool3D_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  maxPool3D_CP_2619_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "maxPool3D_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= maxPool3D_CP_2619_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= maxPool3D_CP_2619_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= maxPool3D_CP_2619_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  maxPool3D_CP_2619: Block -- control-path 
    signal maxPool3D_CP_2619_elements: BooleanArray(202 downto 0);
    -- 
  begin -- 
    maxPool3D_CP_2619_elements(0) <= maxPool3D_CP_2619_start;
    maxPool3D_CP_2619_symbol <= maxPool3D_CP_2619_elements(195);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	37 
    -- CP-element group 0: 	41 
    -- CP-element group 0: 	45 
    -- CP-element group 0: 	49 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	9 
    -- CP-element group 0: 	13 
    -- CP-element group 0: 	17 
    -- CP-element group 0: 	21 
    -- CP-element group 0: 	25 
    -- CP-element group 0: 	29 
    -- CP-element group 0: 	33 
    -- CP-element group 0:  members (44) 
      -- CP-element group 0: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1329_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1346_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1346_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1329_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477__entry__
      -- CP-element group 0: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1358_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1408_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1329_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1396_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1396_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/$entry
      -- CP-element group 0: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1358_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1333_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1371_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1371_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1383_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1333_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1327/$entry
      -- CP-element group 0: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1358_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1383_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1383_Update/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1333_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1346_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1371_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1396_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1408_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1408_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1327/branch_block_stmt_1327__entry__
      -- CP-element group 0: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1421_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1421_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1421_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1433_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1433_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1433_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1446_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1446_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1446_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1458_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1458_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1458_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1471_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1471_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1471_Update/cr
      -- 
    cr_2724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(0), ack => type_cast_1346_inst_req_1); -- 
    cr_2752_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2752_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(0), ack => type_cast_1358_inst_req_1); -- 
    rr_2677_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2677_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(0), ack => RPIPE_maxpool_input_pipe_1329_inst_req_0); -- 
    cr_2836_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2836_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(0), ack => type_cast_1396_inst_req_1); -- 
    cr_2696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(0), ack => type_cast_1333_inst_req_1); -- 
    cr_2780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(0), ack => type_cast_1371_inst_req_1); -- 
    cr_2808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(0), ack => type_cast_1383_inst_req_1); -- 
    cr_2864_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2864_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(0), ack => type_cast_1408_inst_req_1); -- 
    cr_2892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(0), ack => type_cast_1421_inst_req_1); -- 
    cr_2920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(0), ack => type_cast_1433_inst_req_1); -- 
    cr_2948_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2948_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(0), ack => type_cast_1446_inst_req_1); -- 
    cr_2976_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2976_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(0), ack => type_cast_1458_inst_req_1); -- 
    cr_3004_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3004_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(0), ack => type_cast_1471_inst_req_1); -- 
    -- CP-element group 1:  branch  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	182 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	183 
    -- CP-element group 1: 	184 
    -- CP-element group 1:  members (9) 
      -- CP-element group 1: 	 branch_block_stmt_1327/if_stmt_1809_dead_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_1327/if_stmt_1809_eval_test/$entry
      -- CP-element group 1: 	 branch_block_stmt_1327/if_stmt_1809__entry__
      -- CP-element group 1: 	 branch_block_stmt_1327/if_stmt_1809_eval_test/$exit
      -- CP-element group 1: 	 branch_block_stmt_1327/do_while_stmt_1646__exit__
      -- CP-element group 1: 	 branch_block_stmt_1327/if_stmt_1809_else_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_1327/if_stmt_1809_if_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_1327/R_whilex_xbody_whilex_xend_taken_1810_place
      -- CP-element group 1: 	 branch_block_stmt_1327/if_stmt_1809_eval_test/branch_req
      -- 
    branch_req_3455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(1), ack => if_stmt_1809_branch_req_0); -- 
    maxPool3D_CP_2619_elements(1) <= maxPool3D_CP_2619_elements(182);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1329_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1329_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1329_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1329_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1329_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1329_Update/cr
      -- 
    ra_2678_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1329_inst_ack_0, ack => maxPool3D_CP_2619_elements(2)); -- 
    cr_2682_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2682_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(2), ack => RPIPE_maxpool_input_pipe_1329_inst_req_1); -- 
    -- CP-element group 3:  fork  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3: 	6 
    -- CP-element group 3:  members (9) 
      -- CP-element group 3: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1329_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1329_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1329_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1333_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1342_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1342_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1333_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1333_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1342_sample_start_
      -- 
    ca_2683_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1329_inst_ack_1, ack => maxPool3D_CP_2619_elements(3)); -- 
    rr_2691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(3), ack => type_cast_1333_inst_req_0); -- 
    rr_2705_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2705_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(3), ack => RPIPE_maxpool_input_pipe_1342_inst_req_0); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1333_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1333_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1333_sample_completed_
      -- 
    ra_2692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1333_inst_ack_0, ack => maxPool3D_CP_2619_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	50 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1333_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1333_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1333_update_completed_
      -- 
    ca_2697_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1333_inst_ack_1, ack => maxPool3D_CP_2619_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	3 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1342_Update/cr
      -- CP-element group 6: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1342_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1342_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1342_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1342_update_start_
      -- CP-element group 6: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1342_sample_completed_
      -- 
    ra_2706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1342_inst_ack_0, ack => maxPool3D_CP_2619_elements(6)); -- 
    cr_2710_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2710_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(6), ack => RPIPE_maxpool_input_pipe_1342_inst_req_1); -- 
    -- CP-element group 7:  fork  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7: 	10 
    -- CP-element group 7:  members (9) 
      -- CP-element group 7: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1354_Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1342_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1342_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1346_Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1346_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1354_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1342_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1354_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1346_sample_start_
      -- 
    ca_2711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1342_inst_ack_1, ack => maxPool3D_CP_2619_elements(7)); -- 
    rr_2719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(7), ack => type_cast_1346_inst_req_0); -- 
    rr_2733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(7), ack => RPIPE_maxpool_input_pipe_1354_inst_req_0); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1346_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1346_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1346_sample_completed_
      -- 
    ra_2720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1346_inst_ack_0, ack => maxPool3D_CP_2619_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	50 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1346_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1346_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1346_update_completed_
      -- 
    ca_2725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1346_inst_ack_1, ack => maxPool3D_CP_2619_elements(9)); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	7 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1354_update_start_
      -- CP-element group 10: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1354_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1354_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1354_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1354_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1354_Sample/$exit
      -- 
    ra_2734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1354_inst_ack_0, ack => maxPool3D_CP_2619_elements(10)); -- 
    cr_2738_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2738_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(10), ack => RPIPE_maxpool_input_pipe_1354_inst_req_1); -- 
    -- CP-element group 11:  fork  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: 	14 
    -- CP-element group 11:  members (9) 
      -- CP-element group 11: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1354_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1354_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1358_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1367_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1358_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1367_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1358_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1367_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1354_update_completed_
      -- 
    ca_2739_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1354_inst_ack_1, ack => maxPool3D_CP_2619_elements(11)); -- 
    rr_2747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(11), ack => type_cast_1358_inst_req_0); -- 
    rr_2761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(11), ack => RPIPE_maxpool_input_pipe_1367_inst_req_0); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1358_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1358_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1358_sample_completed_
      -- 
    ra_2748_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1358_inst_ack_0, ack => maxPool3D_CP_2619_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	0 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	50 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1358_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1358_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1358_update_completed_
      -- 
    ca_2753_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1358_inst_ack_1, ack => maxPool3D_CP_2619_elements(13)); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	11 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1367_Update/cr
      -- CP-element group 14: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1367_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1367_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1367_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1367_update_start_
      -- CP-element group 14: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1367_sample_completed_
      -- 
    ra_2762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1367_inst_ack_0, ack => maxPool3D_CP_2619_elements(14)); -- 
    cr_2766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(14), ack => RPIPE_maxpool_input_pipe_1367_inst_req_1); -- 
    -- CP-element group 15:  fork  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15: 	18 
    -- CP-element group 15:  members (9) 
      -- CP-element group 15: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1367_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1367_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1379_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1379_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1371_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1371_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1379_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1371_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1367_update_completed_
      -- 
    ca_2767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1367_inst_ack_1, ack => maxPool3D_CP_2619_elements(15)); -- 
    rr_2775_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2775_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(15), ack => type_cast_1371_inst_req_0); -- 
    rr_2789_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2789_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(15), ack => RPIPE_maxpool_input_pipe_1379_inst_req_0); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1371_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1371_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1371_Sample/$exit
      -- 
    ra_2776_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1371_inst_ack_0, ack => maxPool3D_CP_2619_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	0 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	50 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1371_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1371_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1371_update_completed_
      -- 
    ca_2781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1371_inst_ack_1, ack => maxPool3D_CP_2619_elements(17)); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	15 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1379_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1379_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1379_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1379_update_start_
      -- CP-element group 18: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1379_Update/cr
      -- CP-element group 18: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1379_sample_completed_
      -- 
    ra_2790_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1379_inst_ack_0, ack => maxPool3D_CP_2619_elements(18)); -- 
    cr_2794_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2794_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(18), ack => RPIPE_maxpool_input_pipe_1379_inst_req_1); -- 
    -- CP-element group 19:  fork  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19: 	22 
    -- CP-element group 19:  members (9) 
      -- CP-element group 19: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1379_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1383_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1392_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1392_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1383_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1379_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1383_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1392_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1379_Update/$exit
      -- 
    ca_2795_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1379_inst_ack_1, ack => maxPool3D_CP_2619_elements(19)); -- 
    rr_2803_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2803_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(19), ack => type_cast_1383_inst_req_0); -- 
    rr_2817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(19), ack => RPIPE_maxpool_input_pipe_1392_inst_req_0); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1383_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1383_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1383_Sample/ra
      -- 
    ra_2804_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1383_inst_ack_0, ack => maxPool3D_CP_2619_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	0 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	50 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1383_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1383_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1383_Update/$exit
      -- 
    ca_2809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1383_inst_ack_1, ack => maxPool3D_CP_2619_elements(21)); -- 
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	19 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (6) 
      -- CP-element group 22: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1392_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1392_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1392_Update/cr
      -- CP-element group 22: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1392_update_start_
      -- CP-element group 22: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1392_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1392_sample_completed_
      -- 
    ra_2818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1392_inst_ack_0, ack => maxPool3D_CP_2619_elements(22)); -- 
    cr_2822_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2822_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(22), ack => RPIPE_maxpool_input_pipe_1392_inst_req_1); -- 
    -- CP-element group 23:  fork  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: 	26 
    -- CP-element group 23:  members (9) 
      -- CP-element group 23: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1396_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1392_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1404_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1396_Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1404_Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1392_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1404_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1392_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1396_sample_start_
      -- 
    ca_2823_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1392_inst_ack_1, ack => maxPool3D_CP_2619_elements(23)); -- 
    rr_2831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(23), ack => type_cast_1396_inst_req_0); -- 
    rr_2845_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2845_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(23), ack => RPIPE_maxpool_input_pipe_1404_inst_req_0); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1396_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1396_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1396_Sample/ra
      -- 
    ra_2832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1396_inst_ack_0, ack => maxPool3D_CP_2619_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	0 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	50 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1396_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1396_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1396_update_completed_
      -- 
    ca_2837_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1396_inst_ack_1, ack => maxPool3D_CP_2619_elements(25)); -- 
    -- CP-element group 26:  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	23 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (6) 
      -- CP-element group 26: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1404_Update/cr
      -- CP-element group 26: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1404_Update/$entry
      -- CP-element group 26: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1404_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1404_update_start_
      -- CP-element group 26: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1404_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1404_Sample/ra
      -- 
    ra_2846_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1404_inst_ack_0, ack => maxPool3D_CP_2619_elements(26)); -- 
    cr_2850_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2850_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(26), ack => RPIPE_maxpool_input_pipe_1404_inst_req_1); -- 
    -- CP-element group 27:  fork  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27: 	30 
    -- CP-element group 27:  members (9) 
      -- CP-element group 27: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1404_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1417_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1417_Sample/rr
      -- CP-element group 27: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1417_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1404_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1408_Sample/rr
      -- CP-element group 27: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1408_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1408_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1404_Update/$exit
      -- 
    ca_2851_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1404_inst_ack_1, ack => maxPool3D_CP_2619_elements(27)); -- 
    rr_2859_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2859_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(27), ack => type_cast_1408_inst_req_0); -- 
    rr_2873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(27), ack => RPIPE_maxpool_input_pipe_1417_inst_req_0); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1408_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1408_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1408_sample_completed_
      -- 
    ra_2860_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1408_inst_ack_0, ack => maxPool3D_CP_2619_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	0 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	50 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1408_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1408_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1408_Update/ca
      -- 
    ca_2865_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1408_inst_ack_1, ack => maxPool3D_CP_2619_elements(29)); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	27 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1417_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1417_update_start_
      -- CP-element group 30: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1417_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1417_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1417_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1417_Update/cr
      -- 
    ra_2874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1417_inst_ack_0, ack => maxPool3D_CP_2619_elements(30)); -- 
    cr_2878_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2878_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(30), ack => RPIPE_maxpool_input_pipe_1417_inst_req_1); -- 
    -- CP-element group 31:  fork  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31: 	34 
    -- CP-element group 31:  members (9) 
      -- CP-element group 31: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1417_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1417_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1417_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1421_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1421_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1421_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1429_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1429_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1429_Sample/rr
      -- 
    ca_2879_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1417_inst_ack_1, ack => maxPool3D_CP_2619_elements(31)); -- 
    rr_2887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(31), ack => type_cast_1421_inst_req_0); -- 
    rr_2901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(31), ack => RPIPE_maxpool_input_pipe_1429_inst_req_0); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1421_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1421_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1421_Sample/ra
      -- 
    ra_2888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1421_inst_ack_0, ack => maxPool3D_CP_2619_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	0 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	50 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1421_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1421_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1421_Update/ca
      -- 
    ca_2893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1421_inst_ack_1, ack => maxPool3D_CP_2619_elements(33)); -- 
    -- CP-element group 34:  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	31 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (6) 
      -- CP-element group 34: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1429_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1429_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1429_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1429_Sample/ra
      -- CP-element group 34: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1429_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1429_Update/cr
      -- 
    ra_2902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1429_inst_ack_0, ack => maxPool3D_CP_2619_elements(34)); -- 
    cr_2906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(34), ack => RPIPE_maxpool_input_pipe_1429_inst_req_1); -- 
    -- CP-element group 35:  fork  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35: 	38 
    -- CP-element group 35:  members (9) 
      -- CP-element group 35: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1429_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1429_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1429_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1433_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1433_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1433_Sample/rr
      -- CP-element group 35: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1442_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1442_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1442_Sample/rr
      -- 
    ca_2907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1429_inst_ack_1, ack => maxPool3D_CP_2619_elements(35)); -- 
    rr_2929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(35), ack => RPIPE_maxpool_input_pipe_1442_inst_req_0); -- 
    rr_2915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(35), ack => type_cast_1433_inst_req_0); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1433_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1433_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1433_Sample/ra
      -- 
    ra_2916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1433_inst_ack_0, ack => maxPool3D_CP_2619_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	0 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	50 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1433_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1433_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1433_Update/ca
      -- 
    ca_2921_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1433_inst_ack_1, ack => maxPool3D_CP_2619_elements(37)); -- 
    -- CP-element group 38:  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	35 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1442_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1442_update_start_
      -- CP-element group 38: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1442_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1442_Sample/ra
      -- CP-element group 38: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1442_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1442_Update/cr
      -- 
    ra_2930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1442_inst_ack_0, ack => maxPool3D_CP_2619_elements(38)); -- 
    cr_2934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(38), ack => RPIPE_maxpool_input_pipe_1442_inst_req_1); -- 
    -- CP-element group 39:  fork  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39: 	42 
    -- CP-element group 39:  members (9) 
      -- CP-element group 39: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1442_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1442_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1442_Update/ca
      -- CP-element group 39: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1446_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1446_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1446_Sample/rr
      -- CP-element group 39: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1454_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1454_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1454_Sample/rr
      -- 
    ca_2935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1442_inst_ack_1, ack => maxPool3D_CP_2619_elements(39)); -- 
    rr_2943_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2943_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(39), ack => type_cast_1446_inst_req_0); -- 
    rr_2957_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2957_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(39), ack => RPIPE_maxpool_input_pipe_1454_inst_req_0); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1446_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1446_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1446_Sample/ra
      -- 
    ra_2944_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1446_inst_ack_0, ack => maxPool3D_CP_2619_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	0 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	50 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1446_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1446_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1446_Update/ca
      -- 
    ca_2949_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1446_inst_ack_1, ack => maxPool3D_CP_2619_elements(41)); -- 
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	39 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (6) 
      -- CP-element group 42: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1454_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1454_update_start_
      -- CP-element group 42: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1454_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1454_Sample/ra
      -- CP-element group 42: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1454_Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1454_Update/cr
      -- 
    ra_2958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1454_inst_ack_0, ack => maxPool3D_CP_2619_elements(42)); -- 
    cr_2962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(42), ack => RPIPE_maxpool_input_pipe_1454_inst_req_1); -- 
    -- CP-element group 43:  fork  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43: 	46 
    -- CP-element group 43:  members (9) 
      -- CP-element group 43: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1454_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1454_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1454_Update/ca
      -- CP-element group 43: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1458_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1458_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1458_Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1467_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1467_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1467_Sample/rr
      -- 
    ca_2963_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1454_inst_ack_1, ack => maxPool3D_CP_2619_elements(43)); -- 
    rr_2971_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2971_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(43), ack => type_cast_1458_inst_req_0); -- 
    rr_2985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(43), ack => RPIPE_maxpool_input_pipe_1467_inst_req_0); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1458_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1458_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1458_Sample/ra
      -- 
    ra_2972_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1458_inst_ack_0, ack => maxPool3D_CP_2619_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	0 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	50 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1458_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1458_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1458_Update/ca
      -- 
    ca_2977_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1458_inst_ack_1, ack => maxPool3D_CP_2619_elements(45)); -- 
    -- CP-element group 46:  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	43 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (6) 
      -- CP-element group 46: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1467_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1467_update_start_
      -- CP-element group 46: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1467_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1467_Sample/ra
      -- CP-element group 46: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1467_Update/$entry
      -- CP-element group 46: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1467_Update/cr
      -- 
    ra_2986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1467_inst_ack_0, ack => maxPool3D_CP_2619_elements(46)); -- 
    cr_2990_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2990_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(46), ack => RPIPE_maxpool_input_pipe_1467_inst_req_1); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (6) 
      -- CP-element group 47: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1467_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1467_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/RPIPE_maxpool_input_pipe_1467_Update/ca
      -- CP-element group 47: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1471_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1471_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1471_Sample/rr
      -- 
    ca_2991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1467_inst_ack_1, ack => maxPool3D_CP_2619_elements(47)); -- 
    rr_2999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(47), ack => type_cast_1471_inst_req_0); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1471_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1471_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1471_Sample/ra
      -- 
    ra_3000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1471_inst_ack_0, ack => maxPool3D_CP_2619_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	0 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1471_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1471_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/type_cast_1471_Update/ca
      -- 
    ca_3005_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1471_inst_ack_1, ack => maxPool3D_CP_2619_elements(49)); -- 
    -- CP-element group 50:  join  fork  transition  place  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	37 
    -- CP-element group 50: 	41 
    -- CP-element group 50: 	45 
    -- CP-element group 50: 	49 
    -- CP-element group 50: 	5 
    -- CP-element group 50: 	9 
    -- CP-element group 50: 	13 
    -- CP-element group 50: 	17 
    -- CP-element group 50: 	21 
    -- CP-element group 50: 	25 
    -- CP-element group 50: 	29 
    -- CP-element group 50: 	33 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (10) 
      -- CP-element group 50: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477__exit__
      -- CP-element group 50: 	 branch_block_stmt_1327/assign_stmt_1482_to_assign_stmt_1498__entry__
      -- CP-element group 50: 	 branch_block_stmt_1327/assign_stmt_1330_to_assign_stmt_1477/$exit
      -- CP-element group 50: 	 branch_block_stmt_1327/assign_stmt_1482_to_assign_stmt_1498/$entry
      -- CP-element group 50: 	 branch_block_stmt_1327/assign_stmt_1482_to_assign_stmt_1498/type_cast_1481_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_1327/assign_stmt_1482_to_assign_stmt_1498/type_cast_1481_update_start_
      -- CP-element group 50: 	 branch_block_stmt_1327/assign_stmt_1482_to_assign_stmt_1498/type_cast_1481_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_1327/assign_stmt_1482_to_assign_stmt_1498/type_cast_1481_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_1327/assign_stmt_1482_to_assign_stmt_1498/type_cast_1481_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_1327/assign_stmt_1482_to_assign_stmt_1498/type_cast_1481_Update/cr
      -- 
    rr_3016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(50), ack => type_cast_1481_inst_req_0); -- 
    cr_3021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(50), ack => type_cast_1481_inst_req_1); -- 
    maxPool3D_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 11) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_markings: IntegerArray(0 to 11)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant place_delays: IntegerArray(0 to 11) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 12); -- 
    begin -- 
      preds <= maxPool3D_CP_2619_elements(37) & maxPool3D_CP_2619_elements(41) & maxPool3D_CP_2619_elements(45) & maxPool3D_CP_2619_elements(49) & maxPool3D_CP_2619_elements(5) & maxPool3D_CP_2619_elements(9) & maxPool3D_CP_2619_elements(13) & maxPool3D_CP_2619_elements(17) & maxPool3D_CP_2619_elements(21) & maxPool3D_CP_2619_elements(25) & maxPool3D_CP_2619_elements(29) & maxPool3D_CP_2619_elements(33);
      gj_maxPool3D_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 12, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2619_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_1327/assign_stmt_1482_to_assign_stmt_1498/type_cast_1481_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_1327/assign_stmt_1482_to_assign_stmt_1498/type_cast_1481_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_1327/assign_stmt_1482_to_assign_stmt_1498/type_cast_1481_Sample/ra
      -- 
    ra_3017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1481_inst_ack_0, ack => maxPool3D_CP_2619_elements(51)); -- 
    -- CP-element group 52:  branch  transition  place  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (13) 
      -- CP-element group 52: 	 branch_block_stmt_1327/assign_stmt_1482_to_assign_stmt_1498__exit__
      -- CP-element group 52: 	 branch_block_stmt_1327/if_stmt_1499__entry__
      -- CP-element group 52: 	 branch_block_stmt_1327/assign_stmt_1482_to_assign_stmt_1498/$exit
      -- CP-element group 52: 	 branch_block_stmt_1327/assign_stmt_1482_to_assign_stmt_1498/type_cast_1481_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_1327/assign_stmt_1482_to_assign_stmt_1498/type_cast_1481_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_1327/assign_stmt_1482_to_assign_stmt_1498/type_cast_1481_Update/ca
      -- CP-element group 52: 	 branch_block_stmt_1327/if_stmt_1499_dead_link/$entry
      -- CP-element group 52: 	 branch_block_stmt_1327/if_stmt_1499_eval_test/$entry
      -- CP-element group 52: 	 branch_block_stmt_1327/if_stmt_1499_eval_test/$exit
      -- CP-element group 52: 	 branch_block_stmt_1327/if_stmt_1499_eval_test/branch_req
      -- CP-element group 52: 	 branch_block_stmt_1327/R_cmp186_1500_place
      -- CP-element group 52: 	 branch_block_stmt_1327/if_stmt_1499_if_link/$entry
      -- CP-element group 52: 	 branch_block_stmt_1327/if_stmt_1499_else_link/$entry
      -- 
    ca_3022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1481_inst_ack_1, ack => maxPool3D_CP_2619_elements(52)); -- 
    branch_req_3030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(52), ack => if_stmt_1499_branch_req_0); -- 
    -- CP-element group 53:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53: 	56 
    -- CP-element group 53:  members (18) 
      -- CP-element group 53: 	 branch_block_stmt_1327/merge_stmt_1505_PhiAck/$exit
      -- CP-element group 53: 	 branch_block_stmt_1327/assign_stmt_1510_to_assign_stmt_1550__entry__
      -- CP-element group 53: 	 branch_block_stmt_1327/merge_stmt_1505__exit__
      -- CP-element group 53: 	 branch_block_stmt_1327/merge_stmt_1505_PhiAck/$entry
      -- CP-element group 53: 	 branch_block_stmt_1327/merge_stmt_1505_PhiAck/dummy
      -- CP-element group 53: 	 branch_block_stmt_1327/entry_bbx_xnph_PhiReq/$exit
      -- CP-element group 53: 	 branch_block_stmt_1327/entry_bbx_xnph_PhiReq/$entry
      -- CP-element group 53: 	 branch_block_stmt_1327/if_stmt_1499_if_link/$exit
      -- CP-element group 53: 	 branch_block_stmt_1327/if_stmt_1499_if_link/if_choice_transition
      -- CP-element group 53: 	 branch_block_stmt_1327/entry_bbx_xnph
      -- CP-element group 53: 	 branch_block_stmt_1327/merge_stmt_1505_PhiReqMerge
      -- CP-element group 53: 	 branch_block_stmt_1327/assign_stmt_1510_to_assign_stmt_1550/$entry
      -- CP-element group 53: 	 branch_block_stmt_1327/assign_stmt_1510_to_assign_stmt_1550/type_cast_1536_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_1327/assign_stmt_1510_to_assign_stmt_1550/type_cast_1536_update_start_
      -- CP-element group 53: 	 branch_block_stmt_1327/assign_stmt_1510_to_assign_stmt_1550/type_cast_1536_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_1327/assign_stmt_1510_to_assign_stmt_1550/type_cast_1536_Sample/rr
      -- CP-element group 53: 	 branch_block_stmt_1327/assign_stmt_1510_to_assign_stmt_1550/type_cast_1536_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_1327/assign_stmt_1510_to_assign_stmt_1550/type_cast_1536_Update/cr
      -- 
    if_choice_transition_3035_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1499_branch_ack_1, ack => maxPool3D_CP_2619_elements(53)); -- 
    rr_3052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(53), ack => type_cast_1536_inst_req_0); -- 
    cr_3057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(53), ack => type_cast_1536_inst_req_1); -- 
    -- CP-element group 54:  transition  place  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	202 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_1327/if_stmt_1499_else_link/$exit
      -- CP-element group 54: 	 branch_block_stmt_1327/if_stmt_1499_else_link/else_choice_transition
      -- CP-element group 54: 	 branch_block_stmt_1327/entry_forx_xend
      -- CP-element group 54: 	 branch_block_stmt_1327/entry_forx_xend_PhiReq/$entry
      -- CP-element group 54: 	 branch_block_stmt_1327/entry_forx_xend_PhiReq/$exit
      -- 
    else_choice_transition_3039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1499_branch_ack_0, ack => maxPool3D_CP_2619_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_1327/assign_stmt_1510_to_assign_stmt_1550/type_cast_1536_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_1327/assign_stmt_1510_to_assign_stmt_1550/type_cast_1536_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_1327/assign_stmt_1510_to_assign_stmt_1550/type_cast_1536_Sample/ra
      -- 
    ra_3053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1536_inst_ack_0, ack => maxPool3D_CP_2619_elements(55)); -- 
    -- CP-element group 56:  transition  place  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	53 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	196 
    -- CP-element group 56:  members (9) 
      -- CP-element group 56: 	 branch_block_stmt_1327/bbx_xnph_forx_xbody
      -- CP-element group 56: 	 branch_block_stmt_1327/assign_stmt_1510_to_assign_stmt_1550__exit__
      -- CP-element group 56: 	 branch_block_stmt_1327/bbx_xnph_forx_xbody_PhiReq/$entry
      -- CP-element group 56: 	 branch_block_stmt_1327/assign_stmt_1510_to_assign_stmt_1550/$exit
      -- CP-element group 56: 	 branch_block_stmt_1327/assign_stmt_1510_to_assign_stmt_1550/type_cast_1536_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_1327/assign_stmt_1510_to_assign_stmt_1550/type_cast_1536_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_1327/assign_stmt_1510_to_assign_stmt_1550/type_cast_1536_Update/ca
      -- CP-element group 56: 	 branch_block_stmt_1327/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1553/phi_stmt_1553_sources/$entry
      -- CP-element group 56: 	 branch_block_stmt_1327/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1553/$entry
      -- 
    ca_3058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1536_inst_ack_1, ack => maxPool3D_CP_2619_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	201 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_1327/call_stmt_1562_to_assign_stmt_1573/call_stmt_1562_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_1327/call_stmt_1562_to_assign_stmt_1573/call_stmt_1562_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_1327/call_stmt_1562_to_assign_stmt_1573/call_stmt_1562_Sample/cra
      -- 
    cra_3070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1562_call_ack_0, ack => maxPool3D_CP_2619_elements(57)); -- 
    -- CP-element group 58:  branch  transition  place  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	201 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (13) 
      -- CP-element group 58: 	 branch_block_stmt_1327/call_stmt_1562_to_assign_stmt_1573__exit__
      -- CP-element group 58: 	 branch_block_stmt_1327/if_stmt_1574__entry__
      -- CP-element group 58: 	 branch_block_stmt_1327/call_stmt_1562_to_assign_stmt_1573/$exit
      -- CP-element group 58: 	 branch_block_stmt_1327/call_stmt_1562_to_assign_stmt_1573/call_stmt_1562_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_1327/call_stmt_1562_to_assign_stmt_1573/call_stmt_1562_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_1327/call_stmt_1562_to_assign_stmt_1573/call_stmt_1562_Update/cca
      -- CP-element group 58: 	 branch_block_stmt_1327/if_stmt_1574_dead_link/$entry
      -- CP-element group 58: 	 branch_block_stmt_1327/if_stmt_1574_eval_test/$entry
      -- CP-element group 58: 	 branch_block_stmt_1327/if_stmt_1574_eval_test/$exit
      -- CP-element group 58: 	 branch_block_stmt_1327/if_stmt_1574_eval_test/branch_req
      -- CP-element group 58: 	 branch_block_stmt_1327/R_exitcond1_1575_place
      -- CP-element group 58: 	 branch_block_stmt_1327/if_stmt_1574_if_link/$entry
      -- CP-element group 58: 	 branch_block_stmt_1327/if_stmt_1574_else_link/$entry
      -- 
    cca_3075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1562_call_ack_1, ack => maxPool3D_CP_2619_elements(58)); -- 
    branch_req_3083_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3083_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(58), ack => if_stmt_1574_branch_req_0); -- 
    -- CP-element group 59:  merge  transition  place  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	202 
    -- CP-element group 59:  members (13) 
      -- CP-element group 59: 	 branch_block_stmt_1327/merge_stmt_1580_PhiReqMerge
      -- CP-element group 59: 	 branch_block_stmt_1327/merge_stmt_1580__exit__
      -- CP-element group 59: 	 branch_block_stmt_1327/forx_xendx_xloopexit_forx_xend
      -- CP-element group 59: 	 branch_block_stmt_1327/if_stmt_1574_if_link/$exit
      -- CP-element group 59: 	 branch_block_stmt_1327/if_stmt_1574_if_link/if_choice_transition
      -- CP-element group 59: 	 branch_block_stmt_1327/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 59: 	 branch_block_stmt_1327/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_1327/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 59: 	 branch_block_stmt_1327/merge_stmt_1580_PhiAck/$entry
      -- CP-element group 59: 	 branch_block_stmt_1327/merge_stmt_1580_PhiAck/$exit
      -- CP-element group 59: 	 branch_block_stmt_1327/merge_stmt_1580_PhiAck/dummy
      -- CP-element group 59: 	 branch_block_stmt_1327/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_1327/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_3088_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1574_branch_ack_1, ack => maxPool3D_CP_2619_elements(59)); -- 
    -- CP-element group 60:  fork  transition  place  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	197 
    -- CP-element group 60: 	198 
    -- CP-element group 60:  members (12) 
      -- CP-element group 60: 	 branch_block_stmt_1327/forx_xbody_forx_xbody_PhiReq/phi_stmt_1553/phi_stmt_1553_sources/type_cast_1559/SplitProtocol/Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_1327/forx_xbody_forx_xbody_PhiReq/phi_stmt_1553/phi_stmt_1553_sources/type_cast_1559/SplitProtocol/Update/cr
      -- CP-element group 60: 	 branch_block_stmt_1327/forx_xbody_forx_xbody_PhiReq/phi_stmt_1553/phi_stmt_1553_sources/type_cast_1559/SplitProtocol/Sample/rr
      -- CP-element group 60: 	 branch_block_stmt_1327/forx_xbody_forx_xbody_PhiReq/phi_stmt_1553/phi_stmt_1553_sources/type_cast_1559/SplitProtocol/$entry
      -- CP-element group 60: 	 branch_block_stmt_1327/forx_xbody_forx_xbody_PhiReq/phi_stmt_1553/phi_stmt_1553_sources/type_cast_1559/SplitProtocol/Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_1327/forx_xbody_forx_xbody_PhiReq/phi_stmt_1553/phi_stmt_1553_sources/type_cast_1559/$entry
      -- CP-element group 60: 	 branch_block_stmt_1327/forx_xbody_forx_xbody_PhiReq/phi_stmt_1553/phi_stmt_1553_sources/$entry
      -- CP-element group 60: 	 branch_block_stmt_1327/forx_xbody_forx_xbody_PhiReq/phi_stmt_1553/$entry
      -- CP-element group 60: 	 branch_block_stmt_1327/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 60: 	 branch_block_stmt_1327/if_stmt_1574_else_link/$exit
      -- CP-element group 60: 	 branch_block_stmt_1327/if_stmt_1574_else_link/else_choice_transition
      -- CP-element group 60: 	 branch_block_stmt_1327/forx_xbody_forx_xbody
      -- 
    else_choice_transition_3092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1574_branch_ack_0, ack => maxPool3D_CP_2619_elements(60)); -- 
    cr_3588_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3588_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(60), ack => type_cast_1559_inst_req_1); -- 
    rr_3583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(60), ack => type_cast_1559_inst_req_0); -- 
    -- CP-element group 61:  transition  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	202 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_1327/assign_stmt_1599_to_assign_stmt_1603/WPIPE_maxpool_output_pipe_1596_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1327/assign_stmt_1599_to_assign_stmt_1603/WPIPE_maxpool_output_pipe_1596_update_start_
      -- CP-element group 61: 	 branch_block_stmt_1327/assign_stmt_1599_to_assign_stmt_1603/WPIPE_maxpool_output_pipe_1596_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_1327/assign_stmt_1599_to_assign_stmt_1603/WPIPE_maxpool_output_pipe_1596_Sample/ack
      -- CP-element group 61: 	 branch_block_stmt_1327/assign_stmt_1599_to_assign_stmt_1603/WPIPE_maxpool_output_pipe_1596_Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_1327/assign_stmt_1599_to_assign_stmt_1603/WPIPE_maxpool_output_pipe_1596_Update/req
      -- 
    ack_3109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1596_inst_ack_0, ack => maxPool3D_CP_2619_elements(61)); -- 
    req_3113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(61), ack => WPIPE_maxpool_output_pipe_1596_inst_req_1); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (6) 
      -- CP-element group 62: 	 branch_block_stmt_1327/assign_stmt_1599_to_assign_stmt_1603/WPIPE_maxpool_output_pipe_1596_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1327/assign_stmt_1599_to_assign_stmt_1603/WPIPE_maxpool_output_pipe_1596_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_1327/assign_stmt_1599_to_assign_stmt_1603/WPIPE_maxpool_output_pipe_1596_Update/ack
      -- CP-element group 62: 	 branch_block_stmt_1327/assign_stmt_1599_to_assign_stmt_1603/WPIPE_maxpool_output_pipe_1600_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_1327/assign_stmt_1599_to_assign_stmt_1603/WPIPE_maxpool_output_pipe_1600_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_1327/assign_stmt_1599_to_assign_stmt_1603/WPIPE_maxpool_output_pipe_1600_Sample/req
      -- 
    ack_3114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1596_inst_ack_1, ack => maxPool3D_CP_2619_elements(62)); -- 
    req_3122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(62), ack => WPIPE_maxpool_output_pipe_1600_inst_req_0); -- 
    -- CP-element group 63:  transition  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (6) 
      -- CP-element group 63: 	 branch_block_stmt_1327/assign_stmt_1599_to_assign_stmt_1603/WPIPE_maxpool_output_pipe_1600_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_1327/assign_stmt_1599_to_assign_stmt_1603/WPIPE_maxpool_output_pipe_1600_update_start_
      -- CP-element group 63: 	 branch_block_stmt_1327/assign_stmt_1599_to_assign_stmt_1603/WPIPE_maxpool_output_pipe_1600_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_1327/assign_stmt_1599_to_assign_stmt_1603/WPIPE_maxpool_output_pipe_1600_Sample/ack
      -- CP-element group 63: 	 branch_block_stmt_1327/assign_stmt_1599_to_assign_stmt_1603/WPIPE_maxpool_output_pipe_1600_Update/$entry
      -- CP-element group 63: 	 branch_block_stmt_1327/assign_stmt_1599_to_assign_stmt_1603/WPIPE_maxpool_output_pipe_1600_Update/req
      -- 
    ack_3123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1600_inst_ack_0, ack => maxPool3D_CP_2619_elements(63)); -- 
    req_3127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(63), ack => WPIPE_maxpool_output_pipe_1600_inst_req_1); -- 
    -- CP-element group 64:  fork  transition  place  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64: 	66 
    -- CP-element group 64: 	67 
    -- CP-element group 64: 	68 
    -- CP-element group 64: 	69 
    -- CP-element group 64: 	70 
    -- CP-element group 64:  members (25) 
      -- CP-element group 64: 	 branch_block_stmt_1327/assign_stmt_1599_to_assign_stmt_1603__exit__
      -- CP-element group 64: 	 branch_block_stmt_1327/assign_stmt_1608_to_assign_stmt_1627__entry__
      -- CP-element group 64: 	 branch_block_stmt_1327/assign_stmt_1599_to_assign_stmt_1603/$exit
      -- CP-element group 64: 	 branch_block_stmt_1327/assign_stmt_1599_to_assign_stmt_1603/WPIPE_maxpool_output_pipe_1600_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_1327/assign_stmt_1599_to_assign_stmt_1603/WPIPE_maxpool_output_pipe_1600_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_1327/assign_stmt_1599_to_assign_stmt_1603/WPIPE_maxpool_output_pipe_1600_Update/ack
      -- CP-element group 64: 	 branch_block_stmt_1327/assign_stmt_1608_to_assign_stmt_1627/$entry
      -- CP-element group 64: 	 branch_block_stmt_1327/assign_stmt_1608_to_assign_stmt_1627/type_cast_1607_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_1327/assign_stmt_1608_to_assign_stmt_1627/type_cast_1607_update_start_
      -- CP-element group 64: 	 branch_block_stmt_1327/assign_stmt_1608_to_assign_stmt_1627/type_cast_1607_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_1327/assign_stmt_1608_to_assign_stmt_1627/type_cast_1607_Sample/rr
      -- CP-element group 64: 	 branch_block_stmt_1327/assign_stmt_1608_to_assign_stmt_1627/type_cast_1607_Update/$entry
      -- CP-element group 64: 	 branch_block_stmt_1327/assign_stmt_1608_to_assign_stmt_1627/type_cast_1607_Update/cr
      -- CP-element group 64: 	 branch_block_stmt_1327/assign_stmt_1608_to_assign_stmt_1627/type_cast_1611_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_1327/assign_stmt_1608_to_assign_stmt_1627/type_cast_1611_update_start_
      -- CP-element group 64: 	 branch_block_stmt_1327/assign_stmt_1608_to_assign_stmt_1627/type_cast_1611_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_1327/assign_stmt_1608_to_assign_stmt_1627/type_cast_1611_Sample/rr
      -- CP-element group 64: 	 branch_block_stmt_1327/assign_stmt_1608_to_assign_stmt_1627/type_cast_1611_Update/$entry
      -- CP-element group 64: 	 branch_block_stmt_1327/assign_stmt_1608_to_assign_stmt_1627/type_cast_1611_Update/cr
      -- CP-element group 64: 	 branch_block_stmt_1327/assign_stmt_1608_to_assign_stmt_1627/type_cast_1615_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_1327/assign_stmt_1608_to_assign_stmt_1627/type_cast_1615_update_start_
      -- CP-element group 64: 	 branch_block_stmt_1327/assign_stmt_1608_to_assign_stmt_1627/type_cast_1615_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_1327/assign_stmt_1608_to_assign_stmt_1627/type_cast_1615_Sample/rr
      -- CP-element group 64: 	 branch_block_stmt_1327/assign_stmt_1608_to_assign_stmt_1627/type_cast_1615_Update/$entry
      -- CP-element group 64: 	 branch_block_stmt_1327/assign_stmt_1608_to_assign_stmt_1627/type_cast_1615_Update/cr
      -- 
    ack_3128_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1600_inst_ack_1, ack => maxPool3D_CP_2619_elements(64)); -- 
    rr_3139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(64), ack => type_cast_1607_inst_req_0); -- 
    cr_3144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(64), ack => type_cast_1607_inst_req_1); -- 
    rr_3153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(64), ack => type_cast_1611_inst_req_0); -- 
    cr_3158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(64), ack => type_cast_1611_inst_req_1); -- 
    rr_3167_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3167_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(64), ack => type_cast_1615_inst_req_0); -- 
    cr_3172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(64), ack => type_cast_1615_inst_req_1); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_1327/assign_stmt_1608_to_assign_stmt_1627/type_cast_1607_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_1327/assign_stmt_1608_to_assign_stmt_1627/type_cast_1607_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_1327/assign_stmt_1608_to_assign_stmt_1627/type_cast_1607_Sample/ra
      -- 
    ra_3140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1607_inst_ack_0, ack => maxPool3D_CP_2619_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	71 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_1327/assign_stmt_1608_to_assign_stmt_1627/type_cast_1607_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_1327/assign_stmt_1608_to_assign_stmt_1627/type_cast_1607_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_1327/assign_stmt_1608_to_assign_stmt_1627/type_cast_1607_Update/ca
      -- 
    ca_3145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1607_inst_ack_1, ack => maxPool3D_CP_2619_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	64 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1327/assign_stmt_1608_to_assign_stmt_1627/type_cast_1611_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_1327/assign_stmt_1608_to_assign_stmt_1627/type_cast_1611_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_1327/assign_stmt_1608_to_assign_stmt_1627/type_cast_1611_Sample/ra
      -- 
    ra_3154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1611_inst_ack_0, ack => maxPool3D_CP_2619_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	64 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	71 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_1327/assign_stmt_1608_to_assign_stmt_1627/type_cast_1611_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_1327/assign_stmt_1608_to_assign_stmt_1627/type_cast_1611_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_1327/assign_stmt_1608_to_assign_stmt_1627/type_cast_1611_Update/ca
      -- 
    ca_3159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1611_inst_ack_1, ack => maxPool3D_CP_2619_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	64 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_1327/assign_stmt_1608_to_assign_stmt_1627/type_cast_1615_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_1327/assign_stmt_1608_to_assign_stmt_1627/type_cast_1615_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_1327/assign_stmt_1608_to_assign_stmt_1627/type_cast_1615_Sample/ra
      -- 
    ra_3168_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1615_inst_ack_0, ack => maxPool3D_CP_2619_elements(69)); -- 
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	64 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_1327/assign_stmt_1608_to_assign_stmt_1627/type_cast_1615_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_1327/assign_stmt_1608_to_assign_stmt_1627/type_cast_1615_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_1327/assign_stmt_1608_to_assign_stmt_1627/type_cast_1615_Update/ca
      -- 
    ca_3173_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1615_inst_ack_1, ack => maxPool3D_CP_2619_elements(70)); -- 
    -- CP-element group 71:  join  transition  place  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	66 
    -- CP-element group 71: 	68 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (10) 
      -- CP-element group 71: 	 branch_block_stmt_1327/assign_stmt_1608_to_assign_stmt_1627__exit__
      -- CP-element group 71: 	 branch_block_stmt_1327/forx_xend_whilex_xbody
      -- CP-element group 71: 	 branch_block_stmt_1327/merge_stmt_1629__exit__
      -- CP-element group 71: 	 branch_block_stmt_1327/do_while_stmt_1646__entry__
      -- CP-element group 71: 	 branch_block_stmt_1327/assign_stmt_1608_to_assign_stmt_1627/$exit
      -- CP-element group 71: 	 branch_block_stmt_1327/forx_xend_whilex_xbody_PhiReq/$entry
      -- CP-element group 71: 	 branch_block_stmt_1327/forx_xend_whilex_xbody_PhiReq/$exit
      -- CP-element group 71: 	 branch_block_stmt_1327/merge_stmt_1629_PhiReqMerge
      -- CP-element group 71: 	 branch_block_stmt_1327/merge_stmt_1629_PhiAck/$entry
      -- CP-element group 71: 	 branch_block_stmt_1327/merge_stmt_1629_PhiAck/$exit
      -- 
    maxPool3D_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_2619_elements(66) & maxPool3D_CP_2619_elements(68) & maxPool3D_CP_2619_elements(70);
      gj_maxPool3D_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2619_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  transition  place  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	78 
    -- CP-element group 72:  members (2) 
      -- CP-element group 72: 	 branch_block_stmt_1327/do_while_stmt_1646/$entry
      -- CP-element group 72: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646__entry__
      -- 
    maxPool3D_CP_2619_elements(72) <= maxPool3D_CP_2619_elements(71);
    -- CP-element group 73:  merge  place  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	182 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646__exit__
      -- 
    -- Element group maxPool3D_CP_2619_elements(73) is bound as output of CP function.
    -- CP-element group 74:  merge  place  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	77 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_1327/do_while_stmt_1646/loop_back
      -- 
    -- Element group maxPool3D_CP_2619_elements(74) is bound as output of CP function.
    -- CP-element group 75:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	80 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	180 
    -- CP-element group 75: 	181 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_1327/do_while_stmt_1646/loop_taken/$entry
      -- CP-element group 75: 	 branch_block_stmt_1327/do_while_stmt_1646/loop_exit/$entry
      -- CP-element group 75: 	 branch_block_stmt_1327/do_while_stmt_1646/condition_done
      -- 
    maxPool3D_CP_2619_elements(75) <= maxPool3D_CP_2619_elements(80);
    -- CP-element group 76:  branch  place  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	179 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_1327/do_while_stmt_1646/loop_body_done
      -- 
    maxPool3D_CP_2619_elements(76) <= maxPool3D_CP_2619_elements(179);
    -- CP-element group 77:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	74 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	89 
    -- CP-element group 77: 	110 
    -- CP-element group 77: 	131 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/back_edge_to_loop_body
      -- 
    maxPool3D_CP_2619_elements(77) <= maxPool3D_CP_2619_elements(74);
    -- CP-element group 78:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	72 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	91 
    -- CP-element group 78: 	112 
    -- CP-element group 78: 	133 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/first_time_through_loop_body
      -- 
    maxPool3D_CP_2619_elements(78) <= maxPool3D_CP_2619_elements(72);
    -- CP-element group 79:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	85 
    -- CP-element group 79: 	86 
    -- CP-element group 79: 	104 
    -- CP-element group 79: 	105 
    -- CP-element group 79: 	125 
    -- CP-element group 79: 	126 
    -- CP-element group 79: 	178 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/$entry
      -- CP-element group 79: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/loop_body_start
      -- 
    -- Element group maxPool3D_CP_2619_elements(79) is bound as output of CP function.
    -- CP-element group 80:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	84 
    -- CP-element group 80: 	173 
    -- CP-element group 80: 	177 
    -- CP-element group 80: 	178 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	75 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/condition_evaluated
      -- 
    condition_evaluated_3188_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_3188_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(80), ack => do_while_stmt_1646_branch_req_0); -- 
    maxPool3D_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 15);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_2619_elements(84) & maxPool3D_CP_2619_elements(173) & maxPool3D_CP_2619_elements(177) & maxPool3D_CP_2619_elements(178);
      gj_maxPool3D_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2619_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	85 
    -- CP-element group 81: 	104 
    -- CP-element group 81: 	125 
    -- CP-element group 81: marked-predecessors 
    -- CP-element group 81: 	84 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	106 
    -- CP-element group 81: 	127 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/aggregated_phi_sample_req
      -- CP-element group 81: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1648_sample_start__ps
      -- 
    maxPool3D_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_2619_elements(85) & maxPool3D_CP_2619_elements(104) & maxPool3D_CP_2619_elements(125) & maxPool3D_CP_2619_elements(84);
      gj_maxPool3D_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2619_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	87 
    -- CP-element group 82: 	107 
    -- CP-element group 82: 	128 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	163 
    -- CP-element group 82: 	167 
    -- CP-element group 82: 	171 
    -- CP-element group 82: 	175 
    -- CP-element group 82: 	179 
    -- CP-element group 82: marked-successors 
    -- CP-element group 82: 	85 
    -- CP-element group 82: 	104 
    -- CP-element group 82: 	125 
    -- CP-element group 82:  members (4) 
      -- CP-element group 82: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1658_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/aggregated_phi_sample_ack
      -- CP-element group 82: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1648_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1653_sample_completed_
      -- 
    maxPool3D_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_2619_elements(87) & maxPool3D_CP_2619_elements(107) & maxPool3D_CP_2619_elements(128);
      gj_maxPool3D_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2619_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	86 
    -- CP-element group 83: 	105 
    -- CP-element group 83: 	126 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	108 
    -- CP-element group 83: 	129 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/aggregated_phi_update_req
      -- CP-element group 83: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1648_update_start__ps
      -- 
    maxPool3D_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_2619_elements(86) & maxPool3D_CP_2619_elements(105) & maxPool3D_CP_2619_elements(126);
      gj_maxPool3D_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2619_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	88 
    -- CP-element group 84: 	109 
    -- CP-element group 84: 	130 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	80 
    -- CP-element group 84: marked-successors 
    -- CP-element group 84: 	81 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/aggregated_phi_update_ack
      -- 
    maxPool3D_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_2619_elements(88) & maxPool3D_CP_2619_elements(109) & maxPool3D_CP_2619_elements(130);
      gj_maxPool3D_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2619_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  join  transition  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	79 
    -- CP-element group 85: marked-predecessors 
    -- CP-element group 85: 	82 
    -- CP-element group 85: 	173 
    -- CP-element group 85: 	177 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	81 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1648_sample_start_
      -- 
    maxPool3D_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 1,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_2619_elements(79) & maxPool3D_CP_2619_elements(82) & maxPool3D_CP_2619_elements(173) & maxPool3D_CP_2619_elements(177);
      gj_maxPool3D_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2619_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  join  transition  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	79 
    -- CP-element group 86: marked-predecessors 
    -- CP-element group 86: 	88 
    -- CP-element group 86: 	156 
    -- CP-element group 86: 	176 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	83 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1648_update_start_
      -- 
    maxPool3D_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_2619_elements(79) & maxPool3D_CP_2619_elements(88) & maxPool3D_CP_2619_elements(156) & maxPool3D_CP_2619_elements(176);
      gj_maxPool3D_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2619_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  join  transition  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	82 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1648_sample_completed__ps
      -- 
    -- Element group maxPool3D_CP_2619_elements(87) is bound as output of CP function.
    -- CP-element group 88:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	84 
    -- CP-element group 88: 	154 
    -- CP-element group 88: 	174 
    -- CP-element group 88: marked-successors 
    -- CP-element group 88: 	86 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1648_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1648_update_completed__ps
      -- 
    -- Element group maxPool3D_CP_2619_elements(88) is bound as output of CP function.
    -- CP-element group 89:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	77 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (1) 
      -- CP-element group 89: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1648_loopback_trigger
      -- 
    maxPool3D_CP_2619_elements(89) <= maxPool3D_CP_2619_elements(77);
    -- CP-element group 90:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: successors 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1648_loopback_sample_req
      -- CP-element group 90: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1648_loopback_sample_req_ps
      -- 
    phi_stmt_1648_loopback_sample_req_3203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1648_loopback_sample_req_3203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(90), ack => phi_stmt_1648_req_0); -- 
    -- Element group maxPool3D_CP_2619_elements(90) is bound as output of CP function.
    -- CP-element group 91:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	78 
    -- CP-element group 91: successors 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1648_entry_trigger
      -- 
    maxPool3D_CP_2619_elements(91) <= maxPool3D_CP_2619_elements(78);
    -- CP-element group 92:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1648_entry_sample_req
      -- CP-element group 92: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1648_entry_sample_req_ps
      -- 
    phi_stmt_1648_entry_sample_req_3206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1648_entry_sample_req_3206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(92), ack => phi_stmt_1648_req_1); -- 
    -- Element group maxPool3D_CP_2619_elements(92) is bound as output of CP function.
    -- CP-element group 93:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: successors 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1648_phi_mux_ack
      -- CP-element group 93: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1648_phi_mux_ack_ps
      -- 
    phi_stmt_1648_phi_mux_ack_3209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1648_ack_0, ack => maxPool3D_CP_2619_elements(93)); -- 
    -- CP-element group 94:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (1) 
      -- CP-element group 94: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1651_sample_start__ps
      -- 
    -- Element group maxPool3D_CP_2619_elements(94) is bound as output of CP function.
    -- CP-element group 95:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (1) 
      -- CP-element group 95: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1651_update_start__ps
      -- 
    -- Element group maxPool3D_CP_2619_elements(95) is bound as output of CP function.
    -- CP-element group 96:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: marked-predecessors 
    -- CP-element group 96: 	98 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	98 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1651_sample_start_
      -- CP-element group 96: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1651_Sample/$entry
      -- CP-element group 96: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1651_Sample/rr
      -- 
    rr_3222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(96), ack => type_cast_1651_inst_req_0); -- 
    maxPool3D_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2619_elements(94) & maxPool3D_CP_2619_elements(98);
      gj_maxPool3D_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2619_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: marked-predecessors 
    -- CP-element group 97: 	99 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	99 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1651_update_start_
      -- CP-element group 97: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1651_Update/$entry
      -- CP-element group 97: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1651_Update/cr
      -- 
    cr_3227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(97), ack => type_cast_1651_inst_req_1); -- 
    maxPool3D_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2619_elements(95) & maxPool3D_CP_2619_elements(99);
      gj_maxPool3D_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2619_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	96 
    -- CP-element group 98: successors 
    -- CP-element group 98: marked-successors 
    -- CP-element group 98: 	96 
    -- CP-element group 98:  members (4) 
      -- CP-element group 98: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1651_sample_completed__ps
      -- CP-element group 98: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1651_sample_completed_
      -- CP-element group 98: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1651_Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1651_Sample/ra
      -- 
    ra_3223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1651_inst_ack_0, ack => maxPool3D_CP_2619_elements(98)); -- 
    -- CP-element group 99:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	97 
    -- CP-element group 99: successors 
    -- CP-element group 99: marked-successors 
    -- CP-element group 99: 	97 
    -- CP-element group 99:  members (4) 
      -- CP-element group 99: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1651_update_completed__ps
      -- CP-element group 99: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1651_update_completed_
      -- CP-element group 99: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1651_Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1651_Update/ca
      -- 
    ca_3228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1651_inst_ack_1, ack => maxPool3D_CP_2619_elements(99)); -- 
    -- CP-element group 100:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (4) 
      -- CP-element group 100: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/R_rowx_x1_at_entry_1652_sample_start__ps
      -- CP-element group 100: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/R_rowx_x1_at_entry_1652_sample_completed__ps
      -- CP-element group 100: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/R_rowx_x1_at_entry_1652_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/R_rowx_x1_at_entry_1652_sample_completed_
      -- 
    -- Element group maxPool3D_CP_2619_elements(100) is bound as output of CP function.
    -- CP-element group 101:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	103 
    -- CP-element group 101:  members (2) 
      -- CP-element group 101: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/R_rowx_x1_at_entry_1652_update_start__ps
      -- CP-element group 101: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/R_rowx_x1_at_entry_1652_update_start_
      -- 
    -- Element group maxPool3D_CP_2619_elements(101) is bound as output of CP function.
    -- CP-element group 102:  join  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	103 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/R_rowx_x1_at_entry_1652_update_completed__ps
      -- 
    maxPool3D_CP_2619_elements(102) <= maxPool3D_CP_2619_elements(103);
    -- CP-element group 103:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	102 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/R_rowx_x1_at_entry_1652_update_completed_
      -- 
    -- Element group maxPool3D_CP_2619_elements(103) is a control-delay.
    cp_element_103_delay: control_delay_element  generic map(name => " 103_delay", delay_value => 1)  port map(req => maxPool3D_CP_2619_elements(101), ack => maxPool3D_CP_2619_elements(103), clk => clk, reset =>reset);
    -- CP-element group 104:  join  transition  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	79 
    -- CP-element group 104: marked-predecessors 
    -- CP-element group 104: 	82 
    -- CP-element group 104: 	165 
    -- CP-element group 104: 	169 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	81 
    -- CP-element group 104:  members (1) 
      -- CP-element group 104: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1653_sample_start_
      -- 
    maxPool3D_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 1,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_2619_elements(79) & maxPool3D_CP_2619_elements(82) & maxPool3D_CP_2619_elements(165) & maxPool3D_CP_2619_elements(169);
      gj_maxPool3D_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2619_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  join  transition  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	79 
    -- CP-element group 105: marked-predecessors 
    -- CP-element group 105: 	109 
    -- CP-element group 105: 	152 
    -- CP-element group 105: 	168 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	83 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1653_update_start_
      -- 
    maxPool3D_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_2619_elements(79) & maxPool3D_CP_2619_elements(109) & maxPool3D_CP_2619_elements(152) & maxPool3D_CP_2619_elements(168);
      gj_maxPool3D_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2619_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	81 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (1) 
      -- CP-element group 106: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1653_sample_start__ps
      -- 
    maxPool3D_CP_2619_elements(106) <= maxPool3D_CP_2619_elements(81);
    -- CP-element group 107:  join  transition  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	82 
    -- CP-element group 107:  members (1) 
      -- CP-element group 107: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1653_sample_completed__ps
      -- 
    -- Element group maxPool3D_CP_2619_elements(107) is bound as output of CP function.
    -- CP-element group 108:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	83 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1653_update_start__ps
      -- 
    maxPool3D_CP_2619_elements(108) <= maxPool3D_CP_2619_elements(83);
    -- CP-element group 109:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	84 
    -- CP-element group 109: 	150 
    -- CP-element group 109: 	166 
    -- CP-element group 109: marked-successors 
    -- CP-element group 109: 	105 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1653_update_completed_
      -- CP-element group 109: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1653_update_completed__ps
      -- 
    -- Element group maxPool3D_CP_2619_elements(109) is bound as output of CP function.
    -- CP-element group 110:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	77 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1653_loopback_trigger
      -- 
    maxPool3D_CP_2619_elements(110) <= maxPool3D_CP_2619_elements(77);
    -- CP-element group 111:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: successors 
    -- CP-element group 111:  members (2) 
      -- CP-element group 111: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1653_loopback_sample_req
      -- CP-element group 111: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1653_loopback_sample_req_ps
      -- 
    phi_stmt_1653_loopback_sample_req_3247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1653_loopback_sample_req_3247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(111), ack => phi_stmt_1653_req_0); -- 
    -- Element group maxPool3D_CP_2619_elements(111) is bound as output of CP function.
    -- CP-element group 112:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	78 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1653_entry_trigger
      -- 
    maxPool3D_CP_2619_elements(112) <= maxPool3D_CP_2619_elements(78);
    -- CP-element group 113:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: successors 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1653_entry_sample_req
      -- CP-element group 113: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1653_entry_sample_req_ps
      -- 
    phi_stmt_1653_entry_sample_req_3250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1653_entry_sample_req_3250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(113), ack => phi_stmt_1653_req_1); -- 
    -- Element group maxPool3D_CP_2619_elements(113) is bound as output of CP function.
    -- CP-element group 114:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: successors 
    -- CP-element group 114:  members (2) 
      -- CP-element group 114: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1653_phi_mux_ack
      -- CP-element group 114: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1653_phi_mux_ack_ps
      -- 
    phi_stmt_1653_phi_mux_ack_3253_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1653_ack_0, ack => maxPool3D_CP_2619_elements(114)); -- 
    -- CP-element group 115:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (1) 
      -- CP-element group 115: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1656_sample_start__ps
      -- 
    -- Element group maxPool3D_CP_2619_elements(115) is bound as output of CP function.
    -- CP-element group 116:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (1) 
      -- CP-element group 116: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1656_update_start__ps
      -- 
    -- Element group maxPool3D_CP_2619_elements(116) is bound as output of CP function.
    -- CP-element group 117:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: marked-predecessors 
    -- CP-element group 117: 	119 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	119 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1656_Sample/rr
      -- CP-element group 117: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1656_Sample/$entry
      -- CP-element group 117: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1656_sample_start_
      -- 
    rr_3266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(117), ack => type_cast_1656_inst_req_0); -- 
    maxPool3D_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2619_elements(115) & maxPool3D_CP_2619_elements(119);
      gj_maxPool3D_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2619_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: marked-predecessors 
    -- CP-element group 118: 	120 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	120 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1656_Update/cr
      -- CP-element group 118: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1656_Update/$entry
      -- CP-element group 118: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1656_update_start_
      -- 
    cr_3271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(118), ack => type_cast_1656_inst_req_1); -- 
    maxPool3D_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2619_elements(116) & maxPool3D_CP_2619_elements(120);
      gj_maxPool3D_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2619_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	117 
    -- CP-element group 119: successors 
    -- CP-element group 119: marked-successors 
    -- CP-element group 119: 	117 
    -- CP-element group 119:  members (4) 
      -- CP-element group 119: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1656_Sample/ra
      -- CP-element group 119: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1656_Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1656_sample_completed_
      -- CP-element group 119: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1656_sample_completed__ps
      -- 
    ra_3267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1656_inst_ack_0, ack => maxPool3D_CP_2619_elements(119)); -- 
    -- CP-element group 120:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	118 
    -- CP-element group 120: successors 
    -- CP-element group 120: marked-successors 
    -- CP-element group 120: 	118 
    -- CP-element group 120:  members (4) 
      -- CP-element group 120: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1656_Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1656_Update/ca
      -- CP-element group 120: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1656_update_completed_
      -- CP-element group 120: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1656_update_completed__ps
      -- 
    ca_3272_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1656_inst_ack_1, ack => maxPool3D_CP_2619_elements(120)); -- 
    -- CP-element group 121:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (4) 
      -- CP-element group 121: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/R_colx_x1_at_entry_1657_sample_completed__ps
      -- CP-element group 121: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/R_colx_x1_at_entry_1657_sample_start__ps
      -- CP-element group 121: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/R_colx_x1_at_entry_1657_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/R_colx_x1_at_entry_1657_sample_completed_
      -- 
    -- Element group maxPool3D_CP_2619_elements(121) is bound as output of CP function.
    -- CP-element group 122:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	124 
    -- CP-element group 122:  members (2) 
      -- CP-element group 122: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/R_colx_x1_at_entry_1657_update_start__ps
      -- CP-element group 122: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/R_colx_x1_at_entry_1657_update_start_
      -- 
    -- Element group maxPool3D_CP_2619_elements(122) is bound as output of CP function.
    -- CP-element group 123:  join  transition  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	124 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/R_colx_x1_at_entry_1657_update_completed__ps
      -- 
    maxPool3D_CP_2619_elements(123) <= maxPool3D_CP_2619_elements(124);
    -- CP-element group 124:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	122 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	123 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/R_colx_x1_at_entry_1657_update_completed_
      -- 
    -- Element group maxPool3D_CP_2619_elements(124) is a control-delay.
    cp_element_124_delay: control_delay_element  generic map(name => " 124_delay", delay_value => 1)  port map(req => maxPool3D_CP_2619_elements(122), ack => maxPool3D_CP_2619_elements(124), clk => clk, reset =>reset);
    -- CP-element group 125:  join  transition  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	79 
    -- CP-element group 125: marked-predecessors 
    -- CP-element group 125: 	82 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	81 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1658_sample_start_
      -- 
    maxPool3D_cp_element_group_125: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_125"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2619_elements(79) & maxPool3D_CP_2619_elements(82);
      gj_maxPool3D_cp_element_group_125 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2619_elements(125), clk => clk, reset => reset); --
    end block;
    -- CP-element group 126:  join  transition  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	79 
    -- CP-element group 126: marked-predecessors 
    -- CP-element group 126: 	130 
    -- CP-element group 126: 	148 
    -- CP-element group 126: 	164 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	83 
    -- CP-element group 126:  members (1) 
      -- CP-element group 126: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1658_update_start_
      -- 
    maxPool3D_cp_element_group_126: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_126"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_2619_elements(79) & maxPool3D_CP_2619_elements(130) & maxPool3D_CP_2619_elements(148) & maxPool3D_CP_2619_elements(164);
      gj_maxPool3D_cp_element_group_126 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2619_elements(126), clk => clk, reset => reset); --
    end block;
    -- CP-element group 127:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	81 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (1) 
      -- CP-element group 127: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1658_sample_start__ps
      -- 
    maxPool3D_CP_2619_elements(127) <= maxPool3D_CP_2619_elements(81);
    -- CP-element group 128:  join  transition  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	82 
    -- CP-element group 128:  members (1) 
      -- CP-element group 128: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1658_sample_completed__ps
      -- 
    -- Element group maxPool3D_CP_2619_elements(128) is bound as output of CP function.
    -- CP-element group 129:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	83 
    -- CP-element group 129: successors 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1658_update_start__ps
      -- 
    maxPool3D_CP_2619_elements(129) <= maxPool3D_CP_2619_elements(83);
    -- CP-element group 130:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	84 
    -- CP-element group 130: 	146 
    -- CP-element group 130: 	162 
    -- CP-element group 130: marked-successors 
    -- CP-element group 130: 	126 
    -- CP-element group 130:  members (2) 
      -- CP-element group 130: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1658_update_completed_
      -- CP-element group 130: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1658_update_completed__ps
      -- 
    -- Element group maxPool3D_CP_2619_elements(130) is bound as output of CP function.
    -- CP-element group 131:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	77 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (1) 
      -- CP-element group 131: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1658_loopback_trigger
      -- 
    maxPool3D_CP_2619_elements(131) <= maxPool3D_CP_2619_elements(77);
    -- CP-element group 132:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: successors 
    -- CP-element group 132:  members (2) 
      -- CP-element group 132: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1658_loopback_sample_req_ps
      -- CP-element group 132: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1658_loopback_sample_req
      -- 
    phi_stmt_1658_loopback_sample_req_3291_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1658_loopback_sample_req_3291_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(132), ack => phi_stmt_1658_req_0); -- 
    -- Element group maxPool3D_CP_2619_elements(132) is bound as output of CP function.
    -- CP-element group 133:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	78 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (1) 
      -- CP-element group 133: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1658_entry_trigger
      -- 
    maxPool3D_CP_2619_elements(133) <= maxPool3D_CP_2619_elements(78);
    -- CP-element group 134:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: successors 
    -- CP-element group 134:  members (2) 
      -- CP-element group 134: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1658_entry_sample_req_ps
      -- CP-element group 134: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1658_entry_sample_req
      -- 
    phi_stmt_1658_entry_sample_req_3294_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1658_entry_sample_req_3294_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(134), ack => phi_stmt_1658_req_1); -- 
    -- Element group maxPool3D_CP_2619_elements(134) is bound as output of CP function.
    -- CP-element group 135:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (2) 
      -- CP-element group 135: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1658_phi_mux_ack_ps
      -- CP-element group 135: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/phi_stmt_1658_phi_mux_ack
      -- 
    phi_stmt_1658_phi_mux_ack_3297_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1658_ack_0, ack => maxPool3D_CP_2619_elements(135)); -- 
    -- CP-element group 136:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	138 
    -- CP-element group 136:  members (1) 
      -- CP-element group 136: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1661_sample_start__ps
      -- 
    -- Element group maxPool3D_CP_2619_elements(136) is bound as output of CP function.
    -- CP-element group 137:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	139 
    -- CP-element group 137:  members (1) 
      -- CP-element group 137: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1661_update_start__ps
      -- 
    -- Element group maxPool3D_CP_2619_elements(137) is bound as output of CP function.
    -- CP-element group 138:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	136 
    -- CP-element group 138: marked-predecessors 
    -- CP-element group 138: 	140 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	140 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1661_Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1661_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1661_sample_start_
      -- 
    rr_3310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(138), ack => type_cast_1661_inst_req_0); -- 
    maxPool3D_cp_element_group_138: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_138"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2619_elements(136) & maxPool3D_CP_2619_elements(140);
      gj_maxPool3D_cp_element_group_138 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2619_elements(138), clk => clk, reset => reset); --
    end block;
    -- CP-element group 139:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	137 
    -- CP-element group 139: marked-predecessors 
    -- CP-element group 139: 	141 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	141 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1661_Update/cr
      -- CP-element group 139: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1661_Update/$entry
      -- CP-element group 139: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1661_update_start_
      -- 
    cr_3315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(139), ack => type_cast_1661_inst_req_1); -- 
    maxPool3D_cp_element_group_139: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_139"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2619_elements(137) & maxPool3D_CP_2619_elements(141);
      gj_maxPool3D_cp_element_group_139 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2619_elements(139), clk => clk, reset => reset); --
    end block;
    -- CP-element group 140:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	138 
    -- CP-element group 140: successors 
    -- CP-element group 140: marked-successors 
    -- CP-element group 140: 	138 
    -- CP-element group 140:  members (4) 
      -- CP-element group 140: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1661_Sample/ra
      -- CP-element group 140: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1661_Sample/$exit
      -- CP-element group 140: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1661_sample_completed_
      -- CP-element group 140: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1661_sample_completed__ps
      -- 
    ra_3311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1661_inst_ack_0, ack => maxPool3D_CP_2619_elements(140)); -- 
    -- CP-element group 141:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	139 
    -- CP-element group 141: successors 
    -- CP-element group 141: marked-successors 
    -- CP-element group 141: 	139 
    -- CP-element group 141:  members (4) 
      -- CP-element group 141: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1661_Update/ca
      -- CP-element group 141: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1661_Update/$exit
      -- CP-element group 141: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1661_update_completed_
      -- CP-element group 141: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1661_update_completed__ps
      -- 
    ca_3316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1661_inst_ack_1, ack => maxPool3D_CP_2619_elements(141)); -- 
    -- CP-element group 142:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (4) 
      -- CP-element group 142: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/R_chlx_x0_at_entry_1662_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/R_chlx_x0_at_entry_1662_sample_completed__ps
      -- CP-element group 142: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/R_chlx_x0_at_entry_1662_sample_start__ps
      -- CP-element group 142: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/R_chlx_x0_at_entry_1662_sample_completed_
      -- 
    -- Element group maxPool3D_CP_2619_elements(142) is bound as output of CP function.
    -- CP-element group 143:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	145 
    -- CP-element group 143:  members (2) 
      -- CP-element group 143: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/R_chlx_x0_at_entry_1662_update_start__ps
      -- CP-element group 143: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/R_chlx_x0_at_entry_1662_update_start_
      -- 
    -- Element group maxPool3D_CP_2619_elements(143) is bound as output of CP function.
    -- CP-element group 144:  join  transition  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	145 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (1) 
      -- CP-element group 144: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/R_chlx_x0_at_entry_1662_update_completed__ps
      -- 
    maxPool3D_CP_2619_elements(144) <= maxPool3D_CP_2619_elements(145);
    -- CP-element group 145:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	143 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	144 
    -- CP-element group 145:  members (1) 
      -- CP-element group 145: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/R_chlx_x0_at_entry_1662_update_completed_
      -- 
    -- Element group maxPool3D_CP_2619_elements(145) is a control-delay.
    cp_element_145_delay: control_delay_element  generic map(name => " 145_delay", delay_value => 1)  port map(req => maxPool3D_CP_2619_elements(143), ack => maxPool3D_CP_2619_elements(145), clk => clk, reset =>reset);
    -- CP-element group 146:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	130 
    -- CP-element group 146: marked-predecessors 
    -- CP-element group 146: 	148 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	148 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1666_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1666_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1666_Sample/$entry
      -- 
    rr_3333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(146), ack => type_cast_1666_inst_req_0); -- 
    maxPool3D_cp_element_group_146: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_146"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2619_elements(130) & maxPool3D_CP_2619_elements(148);
      gj_maxPool3D_cp_element_group_146 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2619_elements(146), clk => clk, reset => reset); --
    end block;
    -- CP-element group 147:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: marked-predecessors 
    -- CP-element group 147: 	149 
    -- CP-element group 147: 	160 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1666_Update/cr
      -- CP-element group 147: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1666_Update/$entry
      -- CP-element group 147: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1666_update_start_
      -- 
    cr_3338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(147), ack => type_cast_1666_inst_req_1); -- 
    maxPool3D_cp_element_group_147: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_147"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2619_elements(149) & maxPool3D_CP_2619_elements(160);
      gj_maxPool3D_cp_element_group_147 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2619_elements(147), clk => clk, reset => reset); --
    end block;
    -- CP-element group 148:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	146 
    -- CP-element group 148: successors 
    -- CP-element group 148: marked-successors 
    -- CP-element group 148: 	126 
    -- CP-element group 148: 	146 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1666_sample_completed_
      -- CP-element group 148: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1666_Sample/ra
      -- CP-element group 148: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1666_Sample/$exit
      -- 
    ra_3334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1666_inst_ack_0, ack => maxPool3D_CP_2619_elements(148)); -- 
    -- CP-element group 149:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	158 
    -- CP-element group 149: marked-successors 
    -- CP-element group 149: 	147 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1666_Update/ca
      -- CP-element group 149: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1666_Update/$exit
      -- CP-element group 149: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1666_update_completed_
      -- 
    ca_3339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1666_inst_ack_1, ack => maxPool3D_CP_2619_elements(149)); -- 
    -- CP-element group 150:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	109 
    -- CP-element group 150: marked-predecessors 
    -- CP-element group 150: 	152 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1670_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1670_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1670_sample_start_
      -- 
    rr_3347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(150), ack => type_cast_1670_inst_req_0); -- 
    maxPool3D_cp_element_group_150: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_150"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2619_elements(109) & maxPool3D_CP_2619_elements(152);
      gj_maxPool3D_cp_element_group_150 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2619_elements(150), clk => clk, reset => reset); --
    end block;
    -- CP-element group 151:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: marked-predecessors 
    -- CP-element group 151: 	153 
    -- CP-element group 151: 	160 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1670_Update/cr
      -- CP-element group 151: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1670_Update/$entry
      -- CP-element group 151: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1670_update_start_
      -- 
    cr_3352_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3352_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(151), ack => type_cast_1670_inst_req_1); -- 
    maxPool3D_cp_element_group_151: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_151"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2619_elements(153) & maxPool3D_CP_2619_elements(160);
      gj_maxPool3D_cp_element_group_151 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2619_elements(151), clk => clk, reset => reset); --
    end block;
    -- CP-element group 152:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152: marked-successors 
    -- CP-element group 152: 	105 
    -- CP-element group 152: 	150 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1670_Sample/ra
      -- CP-element group 152: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1670_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1670_sample_completed_
      -- 
    ra_3348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1670_inst_ack_0, ack => maxPool3D_CP_2619_elements(152)); -- 
    -- CP-element group 153:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	158 
    -- CP-element group 153: marked-successors 
    -- CP-element group 153: 	151 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1670_Update/ca
      -- CP-element group 153: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1670_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1670_update_completed_
      -- 
    ca_3353_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1670_inst_ack_1, ack => maxPool3D_CP_2619_elements(153)); -- 
    -- CP-element group 154:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	88 
    -- CP-element group 154: marked-predecessors 
    -- CP-element group 154: 	156 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	156 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1674_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1674_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1674_sample_start_
      -- 
    rr_3361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(154), ack => type_cast_1674_inst_req_0); -- 
    maxPool3D_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2619_elements(88) & maxPool3D_CP_2619_elements(156);
      gj_maxPool3D_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2619_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: marked-predecessors 
    -- CP-element group 155: 	157 
    -- CP-element group 155: 	160 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	157 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1674_Update/cr
      -- CP-element group 155: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1674_Update/$entry
      -- CP-element group 155: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1674_update_start_
      -- 
    cr_3366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(155), ack => type_cast_1674_inst_req_1); -- 
    maxPool3D_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2619_elements(157) & maxPool3D_CP_2619_elements(160);
      gj_maxPool3D_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2619_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	154 
    -- CP-element group 156: successors 
    -- CP-element group 156: marked-successors 
    -- CP-element group 156: 	86 
    -- CP-element group 156: 	154 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1674_Sample/ra
      -- CP-element group 156: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1674_Sample/$exit
      -- CP-element group 156: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1674_sample_completed_
      -- 
    ra_3362_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1674_inst_ack_0, ack => maxPool3D_CP_2619_elements(156)); -- 
    -- CP-element group 157:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	158 
    -- CP-element group 157: marked-successors 
    -- CP-element group 157: 	155 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1674_Update/ca
      -- CP-element group 157: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1674_Update/$exit
      -- CP-element group 157: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1674_update_completed_
      -- 
    ca_3367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1674_inst_ack_1, ack => maxPool3D_CP_2619_elements(157)); -- 
    -- CP-element group 158:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	149 
    -- CP-element group 158: 	153 
    -- CP-element group 158: 	157 
    -- CP-element group 158: marked-predecessors 
    -- CP-element group 158: 	160 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	160 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/call_stmt_1743_Sample/crr
      -- CP-element group 158: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/call_stmt_1743_Sample/$entry
      -- CP-element group 158: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/call_stmt_1743_sample_start_
      -- 
    crr_3375_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3375_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(158), ack => call_stmt_1743_call_req_0); -- 
    maxPool3D_cp_element_group_158: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_158"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_2619_elements(149) & maxPool3D_CP_2619_elements(153) & maxPool3D_CP_2619_elements(157) & maxPool3D_CP_2619_elements(160);
      gj_maxPool3D_cp_element_group_158 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2619_elements(158), clk => clk, reset => reset); --
    end block;
    -- CP-element group 159:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: marked-predecessors 
    -- CP-element group 159: 	161 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	161 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/call_stmt_1743_Update/ccr
      -- CP-element group 159: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/call_stmt_1743_Update/$entry
      -- CP-element group 159: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/call_stmt_1743_update_start_
      -- 
    ccr_3380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(159), ack => call_stmt_1743_call_req_1); -- 
    maxPool3D_cp_element_group_159: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_159"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool3D_CP_2619_elements(161);
      gj_maxPool3D_cp_element_group_159 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2619_elements(159), clk => clk, reset => reset); --
    end block;
    -- CP-element group 160:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	158 
    -- CP-element group 160: successors 
    -- CP-element group 160: marked-successors 
    -- CP-element group 160: 	147 
    -- CP-element group 160: 	151 
    -- CP-element group 160: 	155 
    -- CP-element group 160: 	158 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/call_stmt_1743_sample_completed_
      -- CP-element group 160: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/call_stmt_1743_Sample/cra
      -- CP-element group 160: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/call_stmt_1743_Sample/$exit
      -- 
    cra_3376_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1743_call_ack_0, ack => maxPool3D_CP_2619_elements(160)); -- 
    -- CP-element group 161:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	159 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	179 
    -- CP-element group 161: marked-successors 
    -- CP-element group 161: 	159 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/call_stmt_1743_Update/cca
      -- CP-element group 161: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/call_stmt_1743_Update/$exit
      -- CP-element group 161: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/call_stmt_1743_update_completed_
      -- 
    cca_3381_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1743_call_ack_1, ack => maxPool3D_CP_2619_elements(161)); -- 
    -- CP-element group 162:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	130 
    -- CP-element group 162: marked-predecessors 
    -- CP-element group 162: 	164 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	164 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1757_Sample/$entry
      -- CP-element group 162: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1757_sample_start_
      -- CP-element group 162: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1757_Sample/rr
      -- 
    rr_3389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(162), ack => type_cast_1757_inst_req_0); -- 
    maxPool3D_cp_element_group_162: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_162"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2619_elements(130) & maxPool3D_CP_2619_elements(164);
      gj_maxPool3D_cp_element_group_162 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2619_elements(162), clk => clk, reset => reset); --
    end block;
    -- CP-element group 163:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	82 
    -- CP-element group 163: marked-predecessors 
    -- CP-element group 163: 	165 
    -- CP-element group 163: 	172 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	165 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1757_update_start_
      -- CP-element group 163: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1757_Update/cr
      -- CP-element group 163: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1757_Update/$entry
      -- 
    cr_3394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(163), ack => type_cast_1757_inst_req_1); -- 
    maxPool3D_cp_element_group_163: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_163"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_2619_elements(82) & maxPool3D_CP_2619_elements(165) & maxPool3D_CP_2619_elements(172);
      gj_maxPool3D_cp_element_group_163 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2619_elements(163), clk => clk, reset => reset); --
    end block;
    -- CP-element group 164:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	162 
    -- CP-element group 164: successors 
    -- CP-element group 164: marked-successors 
    -- CP-element group 164: 	126 
    -- CP-element group 164: 	162 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1757_sample_completed_
      -- CP-element group 164: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1757_Sample/ra
      -- CP-element group 164: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1757_Sample/$exit
      -- 
    ra_3390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1757_inst_ack_0, ack => maxPool3D_CP_2619_elements(164)); -- 
    -- CP-element group 165:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	163 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	170 
    -- CP-element group 165: marked-successors 
    -- CP-element group 165: 	104 
    -- CP-element group 165: 	163 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1757_update_completed_
      -- CP-element group 165: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1757_Update/ca
      -- CP-element group 165: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1757_Update/$exit
      -- 
    ca_3395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1757_inst_ack_1, ack => maxPool3D_CP_2619_elements(165)); -- 
    -- CP-element group 166:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	109 
    -- CP-element group 166: marked-predecessors 
    -- CP-element group 166: 	168 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	168 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/assign_stmt_1761_Sample/req
      -- CP-element group 166: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/assign_stmt_1761_Sample/$entry
      -- CP-element group 166: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/assign_stmt_1761_sample_start_
      -- 
    req_3403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(166), ack => W_colx_x1_1749_delayed_1_0_1759_inst_req_0); -- 
    maxPool3D_cp_element_group_166: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_166"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2619_elements(109) & maxPool3D_CP_2619_elements(168);
      gj_maxPool3D_cp_element_group_166 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2619_elements(166), clk => clk, reset => reset); --
    end block;
    -- CP-element group 167:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	82 
    -- CP-element group 167: marked-predecessors 
    -- CP-element group 167: 	169 
    -- CP-element group 167: 	172 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	169 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/assign_stmt_1761_update_start_
      -- CP-element group 167: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/assign_stmt_1761_Update/$entry
      -- CP-element group 167: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/assign_stmt_1761_Update/req
      -- 
    req_3408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(167), ack => W_colx_x1_1749_delayed_1_0_1759_inst_req_1); -- 
    maxPool3D_cp_element_group_167: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_167"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_2619_elements(82) & maxPool3D_CP_2619_elements(169) & maxPool3D_CP_2619_elements(172);
      gj_maxPool3D_cp_element_group_167 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2619_elements(167), clk => clk, reset => reset); --
    end block;
    -- CP-element group 168:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	166 
    -- CP-element group 168: successors 
    -- CP-element group 168: marked-successors 
    -- CP-element group 168: 	105 
    -- CP-element group 168: 	166 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/assign_stmt_1761_Sample/ack
      -- CP-element group 168: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/assign_stmt_1761_Sample/$exit
      -- CP-element group 168: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/assign_stmt_1761_sample_completed_
      -- 
    ack_3404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_colx_x1_1749_delayed_1_0_1759_inst_ack_0, ack => maxPool3D_CP_2619_elements(168)); -- 
    -- CP-element group 169:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	170 
    -- CP-element group 169: marked-successors 
    -- CP-element group 169: 	104 
    -- CP-element group 169: 	167 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/assign_stmt_1761_update_completed_
      -- CP-element group 169: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/assign_stmt_1761_Update/ack
      -- CP-element group 169: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/assign_stmt_1761_Update/$exit
      -- 
    ack_3409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_colx_x1_1749_delayed_1_0_1759_inst_ack_1, ack => maxPool3D_CP_2619_elements(169)); -- 
    -- CP-element group 170:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	165 
    -- CP-element group 170: 	169 
    -- CP-element group 170: marked-predecessors 
    -- CP-element group 170: 	172 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	172 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1781_Sample/rr
      -- CP-element group 170: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1781_Sample/$entry
      -- CP-element group 170: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1781_sample_start_
      -- 
    rr_3417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(170), ack => type_cast_1781_inst_req_0); -- 
    maxPool3D_cp_element_group_170: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_170"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_2619_elements(165) & maxPool3D_CP_2619_elements(169) & maxPool3D_CP_2619_elements(172);
      gj_maxPool3D_cp_element_group_170 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2619_elements(170), clk => clk, reset => reset); --
    end block;
    -- CP-element group 171:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	82 
    -- CP-element group 171: marked-predecessors 
    -- CP-element group 171: 	173 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	173 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1781_Update/cr
      -- CP-element group 171: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1781_Update/$entry
      -- CP-element group 171: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1781_update_start_
      -- 
    cr_3422_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3422_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(171), ack => type_cast_1781_inst_req_1); -- 
    maxPool3D_cp_element_group_171: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_171"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2619_elements(82) & maxPool3D_CP_2619_elements(173);
      gj_maxPool3D_cp_element_group_171 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2619_elements(171), clk => clk, reset => reset); --
    end block;
    -- CP-element group 172:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	170 
    -- CP-element group 172: successors 
    -- CP-element group 172: marked-successors 
    -- CP-element group 172: 	163 
    -- CP-element group 172: 	167 
    -- CP-element group 172: 	170 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1781_Sample/ra
      -- CP-element group 172: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1781_Sample/$exit
      -- CP-element group 172: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1781_sample_completed_
      -- 
    ra_3418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1781_inst_ack_0, ack => maxPool3D_CP_2619_elements(172)); -- 
    -- CP-element group 173:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	171 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	80 
    -- CP-element group 173: marked-successors 
    -- CP-element group 173: 	85 
    -- CP-element group 173: 	171 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1781_Update/ca
      -- CP-element group 173: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1781_Update/$exit
      -- CP-element group 173: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/type_cast_1781_update_completed_
      -- 
    ca_3423_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1781_inst_ack_1, ack => maxPool3D_CP_2619_elements(173)); -- 
    -- CP-element group 174:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	88 
    -- CP-element group 174: marked-predecessors 
    -- CP-element group 174: 	176 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	176 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/assign_stmt_1785_Sample/req
      -- CP-element group 174: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/assign_stmt_1785_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/assign_stmt_1785_sample_start_
      -- 
    req_3431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(174), ack => W_rowx_x1_1770_delayed_2_0_1783_inst_req_0); -- 
    maxPool3D_cp_element_group_174: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_174"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2619_elements(88) & maxPool3D_CP_2619_elements(176);
      gj_maxPool3D_cp_element_group_174 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2619_elements(174), clk => clk, reset => reset); --
    end block;
    -- CP-element group 175:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	82 
    -- CP-element group 175: marked-predecessors 
    -- CP-element group 175: 	177 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	177 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/assign_stmt_1785_Update/req
      -- CP-element group 175: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/assign_stmt_1785_Update/$entry
      -- CP-element group 175: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/assign_stmt_1785_update_start_
      -- 
    req_3436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(175), ack => W_rowx_x1_1770_delayed_2_0_1783_inst_req_1); -- 
    maxPool3D_cp_element_group_175: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_175"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2619_elements(82) & maxPool3D_CP_2619_elements(177);
      gj_maxPool3D_cp_element_group_175 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2619_elements(175), clk => clk, reset => reset); --
    end block;
    -- CP-element group 176:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	174 
    -- CP-element group 176: successors 
    -- CP-element group 176: marked-successors 
    -- CP-element group 176: 	86 
    -- CP-element group 176: 	174 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/assign_stmt_1785_Sample/ack
      -- CP-element group 176: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/assign_stmt_1785_Sample/$exit
      -- CP-element group 176: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/assign_stmt_1785_sample_completed_
      -- 
    ack_3432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rowx_x1_1770_delayed_2_0_1783_inst_ack_0, ack => maxPool3D_CP_2619_elements(176)); -- 
    -- CP-element group 177:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	175 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	80 
    -- CP-element group 177: marked-successors 
    -- CP-element group 177: 	85 
    -- CP-element group 177: 	175 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/assign_stmt_1785_Update/ack
      -- CP-element group 177: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/assign_stmt_1785_Update/$exit
      -- CP-element group 177: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/assign_stmt_1785_update_completed_
      -- 
    ack_3437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rowx_x1_1770_delayed_2_0_1783_inst_ack_1, ack => maxPool3D_CP_2619_elements(177)); -- 
    -- CP-element group 178:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	79 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	80 
    -- CP-element group 178:  members (1) 
      -- CP-element group 178: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group maxPool3D_CP_2619_elements(178) is a control-delay.
    cp_element_178_delay: control_delay_element  generic map(name => " 178_delay", delay_value => 1)  port map(req => maxPool3D_CP_2619_elements(79), ack => maxPool3D_CP_2619_elements(178), clk => clk, reset =>reset);
    -- CP-element group 179:  join  transition  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	82 
    -- CP-element group 179: 	161 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	76 
    -- CP-element group 179:  members (1) 
      -- CP-element group 179: 	 branch_block_stmt_1327/do_while_stmt_1646/do_while_stmt_1646_loop_body/$exit
      -- 
    maxPool3D_cp_element_group_179: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_179"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2619_elements(82) & maxPool3D_CP_2619_elements(161);
      gj_maxPool3D_cp_element_group_179 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2619_elements(179), clk => clk, reset => reset); --
    end block;
    -- CP-element group 180:  transition  input  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	75 
    -- CP-element group 180: successors 
    -- CP-element group 180:  members (2) 
      -- CP-element group 180: 	 branch_block_stmt_1327/do_while_stmt_1646/loop_exit/ack
      -- CP-element group 180: 	 branch_block_stmt_1327/do_while_stmt_1646/loop_exit/$exit
      -- 
    ack_3442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1646_branch_ack_0, ack => maxPool3D_CP_2619_elements(180)); -- 
    -- CP-element group 181:  transition  input  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	75 
    -- CP-element group 181: successors 
    -- CP-element group 181:  members (2) 
      -- CP-element group 181: 	 branch_block_stmt_1327/do_while_stmt_1646/loop_taken/ack
      -- CP-element group 181: 	 branch_block_stmt_1327/do_while_stmt_1646/loop_taken/$exit
      -- 
    ack_3446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1646_branch_ack_1, ack => maxPool3D_CP_2619_elements(181)); -- 
    -- CP-element group 182:  transition  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	73 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	1 
    -- CP-element group 182:  members (1) 
      -- CP-element group 182: 	 branch_block_stmt_1327/do_while_stmt_1646/$exit
      -- 
    maxPool3D_CP_2619_elements(182) <= maxPool3D_CP_2619_elements(73);
    -- CP-element group 183:  merge  transition  place  input  output  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	1 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	185 
    -- CP-element group 183:  members (15) 
      -- CP-element group 183: 	 branch_block_stmt_1327/merge_stmt_1813__exit__
      -- CP-element group 183: 	 branch_block_stmt_1327/assign_stmt_1818_to_assign_stmt_1822/WPIPE_maxpool_output_pipe_1815_Sample/$entry
      -- CP-element group 183: 	 branch_block_stmt_1327/assign_stmt_1818_to_assign_stmt_1822__entry__
      -- CP-element group 183: 	 branch_block_stmt_1327/assign_stmt_1818_to_assign_stmt_1822/WPIPE_maxpool_output_pipe_1815_Sample/req
      -- CP-element group 183: 	 branch_block_stmt_1327/assign_stmt_1818_to_assign_stmt_1822/WPIPE_maxpool_output_pipe_1815_sample_start_
      -- CP-element group 183: 	 branch_block_stmt_1327/assign_stmt_1818_to_assign_stmt_1822/$entry
      -- CP-element group 183: 	 branch_block_stmt_1327/if_stmt_1809_if_link/if_choice_transition
      -- CP-element group 183: 	 branch_block_stmt_1327/if_stmt_1809_if_link/$exit
      -- CP-element group 183: 	 branch_block_stmt_1327/whilex_xbody_whilex_xend
      -- CP-element group 183: 	 branch_block_stmt_1327/whilex_xbody_whilex_xend_PhiReq/$entry
      -- CP-element group 183: 	 branch_block_stmt_1327/whilex_xbody_whilex_xend_PhiReq/$exit
      -- CP-element group 183: 	 branch_block_stmt_1327/merge_stmt_1813_PhiReqMerge
      -- CP-element group 183: 	 branch_block_stmt_1327/merge_stmt_1813_PhiAck/$entry
      -- CP-element group 183: 	 branch_block_stmt_1327/merge_stmt_1813_PhiAck/$exit
      -- CP-element group 183: 	 branch_block_stmt_1327/merge_stmt_1813_PhiAck/dummy
      -- 
    if_choice_transition_3460_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1809_branch_ack_1, ack => maxPool3D_CP_2619_elements(183)); -- 
    req_3476_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3476_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(183), ack => WPIPE_maxpool_output_pipe_1815_inst_req_0); -- 
    -- CP-element group 184:  merge  transition  place  input  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	1 
    -- CP-element group 184: successors 
    -- CP-element group 184:  members (5) 
      -- CP-element group 184: 	 branch_block_stmt_1327/merge_stmt_1813__entry__
      -- CP-element group 184: 	 branch_block_stmt_1327/if_stmt_1809__exit__
      -- CP-element group 184: 	 branch_block_stmt_1327/if_stmt_1809_else_link/else_choice_transition
      -- CP-element group 184: 	 branch_block_stmt_1327/if_stmt_1809_else_link/$exit
      -- CP-element group 184: 	 branch_block_stmt_1327/merge_stmt_1813_dead_link/$entry
      -- 
    else_choice_transition_3464_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1809_branch_ack_0, ack => maxPool3D_CP_2619_elements(184)); -- 
    -- CP-element group 185:  transition  input  output  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	183 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	186 
    -- CP-element group 185:  members (6) 
      -- CP-element group 185: 	 branch_block_stmt_1327/assign_stmt_1818_to_assign_stmt_1822/WPIPE_maxpool_output_pipe_1815_Sample/$exit
      -- CP-element group 185: 	 branch_block_stmt_1327/assign_stmt_1818_to_assign_stmt_1822/WPIPE_maxpool_output_pipe_1815_Update/$entry
      -- CP-element group 185: 	 branch_block_stmt_1327/assign_stmt_1818_to_assign_stmt_1822/WPIPE_maxpool_output_pipe_1815_Update/req
      -- CP-element group 185: 	 branch_block_stmt_1327/assign_stmt_1818_to_assign_stmt_1822/WPIPE_maxpool_output_pipe_1815_Sample/ack
      -- CP-element group 185: 	 branch_block_stmt_1327/assign_stmt_1818_to_assign_stmt_1822/WPIPE_maxpool_output_pipe_1815_update_start_
      -- CP-element group 185: 	 branch_block_stmt_1327/assign_stmt_1818_to_assign_stmt_1822/WPIPE_maxpool_output_pipe_1815_sample_completed_
      -- 
    ack_3477_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1815_inst_ack_0, ack => maxPool3D_CP_2619_elements(185)); -- 
    req_3481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(185), ack => WPIPE_maxpool_output_pipe_1815_inst_req_1); -- 
    -- CP-element group 186:  transition  input  output  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	185 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186:  members (6) 
      -- CP-element group 186: 	 branch_block_stmt_1327/assign_stmt_1818_to_assign_stmt_1822/WPIPE_maxpool_output_pipe_1815_Update/ack
      -- CP-element group 186: 	 branch_block_stmt_1327/assign_stmt_1818_to_assign_stmt_1822/WPIPE_maxpool_output_pipe_1819_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_1327/assign_stmt_1818_to_assign_stmt_1822/WPIPE_maxpool_output_pipe_1819_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_1327/assign_stmt_1818_to_assign_stmt_1822/WPIPE_maxpool_output_pipe_1815_Update/$exit
      -- CP-element group 186: 	 branch_block_stmt_1327/assign_stmt_1818_to_assign_stmt_1822/WPIPE_maxpool_output_pipe_1815_update_completed_
      -- CP-element group 186: 	 branch_block_stmt_1327/assign_stmt_1818_to_assign_stmt_1822/WPIPE_maxpool_output_pipe_1819_Sample/req
      -- 
    ack_3482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1815_inst_ack_1, ack => maxPool3D_CP_2619_elements(186)); -- 
    req_3490_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3490_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(186), ack => WPIPE_maxpool_output_pipe_1819_inst_req_0); -- 
    -- CP-element group 187:  transition  input  output  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187:  members (6) 
      -- CP-element group 187: 	 branch_block_stmt_1327/assign_stmt_1818_to_assign_stmt_1822/WPIPE_maxpool_output_pipe_1819_update_start_
      -- CP-element group 187: 	 branch_block_stmt_1327/assign_stmt_1818_to_assign_stmt_1822/WPIPE_maxpool_output_pipe_1819_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_1327/assign_stmt_1818_to_assign_stmt_1822/WPIPE_maxpool_output_pipe_1819_Sample/$exit
      -- CP-element group 187: 	 branch_block_stmt_1327/assign_stmt_1818_to_assign_stmt_1822/WPIPE_maxpool_output_pipe_1819_Update/req
      -- CP-element group 187: 	 branch_block_stmt_1327/assign_stmt_1818_to_assign_stmt_1822/WPIPE_maxpool_output_pipe_1819_Update/$entry
      -- CP-element group 187: 	 branch_block_stmt_1327/assign_stmt_1818_to_assign_stmt_1822/WPIPE_maxpool_output_pipe_1819_Sample/ack
      -- 
    ack_3491_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1819_inst_ack_0, ack => maxPool3D_CP_2619_elements(187)); -- 
    req_3495_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3495_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(187), ack => WPIPE_maxpool_output_pipe_1819_inst_req_1); -- 
    -- CP-element group 188:  fork  transition  place  input  output  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	189 
    -- CP-element group 188: 	190 
    -- CP-element group 188: 	191 
    -- CP-element group 188: 	192 
    -- CP-element group 188: 	195 
    -- CP-element group 188:  members (22) 
      -- CP-element group 188: 	 branch_block_stmt_1327/assign_stmt_1818_to_assign_stmt_1822/WPIPE_maxpool_output_pipe_1819_update_completed_
      -- CP-element group 188: 	 branch_block_stmt_1327/assign_stmt_1827_to_call_stmt_1843/type_cast_1830_Sample/rr
      -- CP-element group 188: 	 branch_block_stmt_1327/assign_stmt_1827_to_call_stmt_1843/type_cast_1830_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_1327/assign_stmt_1827_to_call_stmt_1843/type_cast_1826_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_1327/assign_stmt_1827_to_call_stmt_1843__entry__
      -- CP-element group 188: 	 branch_block_stmt_1327/assign_stmt_1818_to_assign_stmt_1822__exit__
      -- CP-element group 188: 	 branch_block_stmt_1327/assign_stmt_1827_to_call_stmt_1843/type_cast_1826_Sample/rr
      -- CP-element group 188: 	 branch_block_stmt_1327/assign_stmt_1827_to_call_stmt_1843/type_cast_1826_update_start_
      -- CP-element group 188: 	 branch_block_stmt_1327/assign_stmt_1818_to_assign_stmt_1822/$exit
      -- CP-element group 188: 	 branch_block_stmt_1327/assign_stmt_1827_to_call_stmt_1843/type_cast_1826_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_1327/assign_stmt_1827_to_call_stmt_1843/$entry
      -- CP-element group 188: 	 branch_block_stmt_1327/assign_stmt_1827_to_call_stmt_1843/call_stmt_1843_Update/ccr
      -- CP-element group 188: 	 branch_block_stmt_1327/assign_stmt_1818_to_assign_stmt_1822/WPIPE_maxpool_output_pipe_1819_Update/ack
      -- CP-element group 188: 	 branch_block_stmt_1327/assign_stmt_1818_to_assign_stmt_1822/WPIPE_maxpool_output_pipe_1819_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_1327/assign_stmt_1827_to_call_stmt_1843/call_stmt_1843_Update/$entry
      -- CP-element group 188: 	 branch_block_stmt_1327/assign_stmt_1827_to_call_stmt_1843/type_cast_1830_update_start_
      -- CP-element group 188: 	 branch_block_stmt_1327/assign_stmt_1827_to_call_stmt_1843/type_cast_1830_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_1327/assign_stmt_1827_to_call_stmt_1843/type_cast_1826_Update/cr
      -- CP-element group 188: 	 branch_block_stmt_1327/assign_stmt_1827_to_call_stmt_1843/call_stmt_1843_update_start_
      -- CP-element group 188: 	 branch_block_stmt_1327/assign_stmt_1827_to_call_stmt_1843/type_cast_1826_Update/$entry
      -- CP-element group 188: 	 branch_block_stmt_1327/assign_stmt_1827_to_call_stmt_1843/type_cast_1830_Update/cr
      -- CP-element group 188: 	 branch_block_stmt_1327/assign_stmt_1827_to_call_stmt_1843/type_cast_1830_Update/$entry
      -- 
    ack_3496_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1819_inst_ack_1, ack => maxPool3D_CP_2619_elements(188)); -- 
    rr_3521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(188), ack => type_cast_1830_inst_req_0); -- 
    rr_3507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(188), ack => type_cast_1826_inst_req_0); -- 
    ccr_3540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(188), ack => call_stmt_1843_call_req_1); -- 
    cr_3512_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3512_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(188), ack => type_cast_1826_inst_req_1); -- 
    cr_3526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(188), ack => type_cast_1830_inst_req_1); -- 
    -- CP-element group 189:  transition  input  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	188 
    -- CP-element group 189: successors 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_1327/assign_stmt_1827_to_call_stmt_1843/type_cast_1826_Sample/$exit
      -- CP-element group 189: 	 branch_block_stmt_1327/assign_stmt_1827_to_call_stmt_1843/type_cast_1826_Sample/ra
      -- CP-element group 189: 	 branch_block_stmt_1327/assign_stmt_1827_to_call_stmt_1843/type_cast_1826_sample_completed_
      -- 
    ra_3508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1826_inst_ack_0, ack => maxPool3D_CP_2619_elements(189)); -- 
    -- CP-element group 190:  transition  input  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	188 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	193 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_1327/assign_stmt_1827_to_call_stmt_1843/type_cast_1826_update_completed_
      -- CP-element group 190: 	 branch_block_stmt_1327/assign_stmt_1827_to_call_stmt_1843/type_cast_1826_Update/ca
      -- CP-element group 190: 	 branch_block_stmt_1327/assign_stmt_1827_to_call_stmt_1843/type_cast_1826_Update/$exit
      -- 
    ca_3513_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1826_inst_ack_1, ack => maxPool3D_CP_2619_elements(190)); -- 
    -- CP-element group 191:  transition  input  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	188 
    -- CP-element group 191: successors 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_1327/assign_stmt_1827_to_call_stmt_1843/type_cast_1830_Sample/ra
      -- CP-element group 191: 	 branch_block_stmt_1327/assign_stmt_1827_to_call_stmt_1843/type_cast_1830_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_1327/assign_stmt_1827_to_call_stmt_1843/type_cast_1830_sample_completed_
      -- 
    ra_3522_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1830_inst_ack_0, ack => maxPool3D_CP_2619_elements(191)); -- 
    -- CP-element group 192:  transition  input  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	188 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	193 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_1327/assign_stmt_1827_to_call_stmt_1843/type_cast_1830_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_1327/assign_stmt_1827_to_call_stmt_1843/type_cast_1830_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_1327/assign_stmt_1827_to_call_stmt_1843/type_cast_1830_Update/ca
      -- 
    ca_3527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1830_inst_ack_1, ack => maxPool3D_CP_2619_elements(192)); -- 
    -- CP-element group 193:  join  transition  output  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	190 
    -- CP-element group 193: 	192 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	194 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_1327/assign_stmt_1827_to_call_stmt_1843/call_stmt_1843_Sample/crr
      -- CP-element group 193: 	 branch_block_stmt_1327/assign_stmt_1827_to_call_stmt_1843/call_stmt_1843_Sample/$entry
      -- CP-element group 193: 	 branch_block_stmt_1327/assign_stmt_1827_to_call_stmt_1843/call_stmt_1843_sample_start_
      -- 
    crr_3535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(193), ack => call_stmt_1843_call_req_0); -- 
    maxPool3D_cp_element_group_193: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_193"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2619_elements(190) & maxPool3D_CP_2619_elements(192);
      gj_maxPool3D_cp_element_group_193 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2619_elements(193), clk => clk, reset => reset); --
    end block;
    -- CP-element group 194:  transition  input  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	193 
    -- CP-element group 194: successors 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_1327/assign_stmt_1827_to_call_stmt_1843/call_stmt_1843_Sample/cra
      -- CP-element group 194: 	 branch_block_stmt_1327/assign_stmt_1827_to_call_stmt_1843/call_stmt_1843_Sample/$exit
      -- CP-element group 194: 	 branch_block_stmt_1327/assign_stmt_1827_to_call_stmt_1843/call_stmt_1843_sample_completed_
      -- 
    cra_3536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1843_call_ack_0, ack => maxPool3D_CP_2619_elements(194)); -- 
    -- CP-element group 195:  transition  place  input  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	188 
    -- CP-element group 195: successors 
    -- CP-element group 195:  members (16) 
      -- CP-element group 195: 	 branch_block_stmt_1327/branch_block_stmt_1327__exit__
      -- CP-element group 195: 	 branch_block_stmt_1327/merge_stmt_1845__exit__
      -- CP-element group 195: 	 branch_block_stmt_1327/return__
      -- CP-element group 195: 	 branch_block_stmt_1327/assign_stmt_1827_to_call_stmt_1843__exit__
      -- CP-element group 195: 	 branch_block_stmt_1327/$exit
      -- CP-element group 195: 	 $exit
      -- CP-element group 195: 	 branch_block_stmt_1327/assign_stmt_1827_to_call_stmt_1843/$exit
      -- CP-element group 195: 	 branch_block_stmt_1327/assign_stmt_1827_to_call_stmt_1843/call_stmt_1843_Update/cca
      -- CP-element group 195: 	 branch_block_stmt_1327/assign_stmt_1827_to_call_stmt_1843/call_stmt_1843_Update/$exit
      -- CP-element group 195: 	 branch_block_stmt_1327/assign_stmt_1827_to_call_stmt_1843/call_stmt_1843_update_completed_
      -- CP-element group 195: 	 branch_block_stmt_1327/return___PhiReq/$entry
      -- CP-element group 195: 	 branch_block_stmt_1327/return___PhiReq/$exit
      -- CP-element group 195: 	 branch_block_stmt_1327/merge_stmt_1845_PhiReqMerge
      -- CP-element group 195: 	 branch_block_stmt_1327/merge_stmt_1845_PhiAck/$entry
      -- CP-element group 195: 	 branch_block_stmt_1327/merge_stmt_1845_PhiAck/$exit
      -- CP-element group 195: 	 branch_block_stmt_1327/merge_stmt_1845_PhiAck/dummy
      -- 
    cca_3541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1843_call_ack_1, ack => maxPool3D_CP_2619_elements(195)); -- 
    -- CP-element group 196:  transition  output  delay-element  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	56 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	200 
    -- CP-element group 196:  members (5) 
      -- CP-element group 196: 	 branch_block_stmt_1327/bbx_xnph_forx_xbody_PhiReq/$exit
      -- CP-element group 196: 	 branch_block_stmt_1327/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1553/phi_stmt_1553_req
      -- CP-element group 196: 	 branch_block_stmt_1327/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1553/phi_stmt_1553_sources/type_cast_1557_konst_delay_trans
      -- CP-element group 196: 	 branch_block_stmt_1327/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1553/phi_stmt_1553_sources/$exit
      -- CP-element group 196: 	 branch_block_stmt_1327/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1553/$exit
      -- 
    phi_stmt_1553_req_3564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1553_req_3564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(196), ack => phi_stmt_1553_req_0); -- 
    -- Element group maxPool3D_CP_2619_elements(196) is a control-delay.
    cp_element_196_delay: control_delay_element  generic map(name => " 196_delay", delay_value => 1)  port map(req => maxPool3D_CP_2619_elements(56), ack => maxPool3D_CP_2619_elements(196), clk => clk, reset =>reset);
    -- CP-element group 197:  transition  input  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	60 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	199 
    -- CP-element group 197:  members (2) 
      -- CP-element group 197: 	 branch_block_stmt_1327/forx_xbody_forx_xbody_PhiReq/phi_stmt_1553/phi_stmt_1553_sources/type_cast_1559/SplitProtocol/Sample/ra
      -- CP-element group 197: 	 branch_block_stmt_1327/forx_xbody_forx_xbody_PhiReq/phi_stmt_1553/phi_stmt_1553_sources/type_cast_1559/SplitProtocol/Sample/$exit
      -- 
    ra_3584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1559_inst_ack_0, ack => maxPool3D_CP_2619_elements(197)); -- 
    -- CP-element group 198:  transition  input  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	60 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	199 
    -- CP-element group 198:  members (2) 
      -- CP-element group 198: 	 branch_block_stmt_1327/forx_xbody_forx_xbody_PhiReq/phi_stmt_1553/phi_stmt_1553_sources/type_cast_1559/SplitProtocol/Update/$exit
      -- CP-element group 198: 	 branch_block_stmt_1327/forx_xbody_forx_xbody_PhiReq/phi_stmt_1553/phi_stmt_1553_sources/type_cast_1559/SplitProtocol/Update/ca
      -- 
    ca_3589_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1559_inst_ack_1, ack => maxPool3D_CP_2619_elements(198)); -- 
    -- CP-element group 199:  join  transition  output  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	197 
    -- CP-element group 199: 	198 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199:  members (6) 
      -- CP-element group 199: 	 branch_block_stmt_1327/forx_xbody_forx_xbody_PhiReq/phi_stmt_1553/phi_stmt_1553_req
      -- CP-element group 199: 	 branch_block_stmt_1327/forx_xbody_forx_xbody_PhiReq/phi_stmt_1553/phi_stmt_1553_sources/type_cast_1559/SplitProtocol/$exit
      -- CP-element group 199: 	 branch_block_stmt_1327/forx_xbody_forx_xbody_PhiReq/phi_stmt_1553/phi_stmt_1553_sources/type_cast_1559/$exit
      -- CP-element group 199: 	 branch_block_stmt_1327/forx_xbody_forx_xbody_PhiReq/phi_stmt_1553/phi_stmt_1553_sources/$exit
      -- CP-element group 199: 	 branch_block_stmt_1327/forx_xbody_forx_xbody_PhiReq/phi_stmt_1553/$exit
      -- CP-element group 199: 	 branch_block_stmt_1327/forx_xbody_forx_xbody_PhiReq/$exit
      -- 
    phi_stmt_1553_req_3590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1553_req_3590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(199), ack => phi_stmt_1553_req_1); -- 
    maxPool3D_cp_element_group_199: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_199"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2619_elements(197) & maxPool3D_CP_2619_elements(198);
      gj_maxPool3D_cp_element_group_199 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2619_elements(199), clk => clk, reset => reset); --
    end block;
    -- CP-element group 200:  merge  transition  place  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	196 
    -- CP-element group 200: 	199 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	201 
    -- CP-element group 200:  members (2) 
      -- CP-element group 200: 	 branch_block_stmt_1327/merge_stmt_1552_PhiAck/$entry
      -- CP-element group 200: 	 branch_block_stmt_1327/merge_stmt_1552_PhiReqMerge
      -- 
    maxPool3D_CP_2619_elements(200) <= OrReduce(maxPool3D_CP_2619_elements(196) & maxPool3D_CP_2619_elements(199));
    -- CP-element group 201:  fork  transition  place  input  output  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	200 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	57 
    -- CP-element group 201: 	58 
    -- CP-element group 201:  members (11) 
      -- CP-element group 201: 	 branch_block_stmt_1327/merge_stmt_1552__exit__
      -- CP-element group 201: 	 branch_block_stmt_1327/call_stmt_1562_to_assign_stmt_1573__entry__
      -- CP-element group 201: 	 branch_block_stmt_1327/merge_stmt_1552_PhiAck/$exit
      -- CP-element group 201: 	 branch_block_stmt_1327/merge_stmt_1552_PhiAck/phi_stmt_1553_ack
      -- CP-element group 201: 	 branch_block_stmt_1327/call_stmt_1562_to_assign_stmt_1573/$entry
      -- CP-element group 201: 	 branch_block_stmt_1327/call_stmt_1562_to_assign_stmt_1573/call_stmt_1562_sample_start_
      -- CP-element group 201: 	 branch_block_stmt_1327/call_stmt_1562_to_assign_stmt_1573/call_stmt_1562_update_start_
      -- CP-element group 201: 	 branch_block_stmt_1327/call_stmt_1562_to_assign_stmt_1573/call_stmt_1562_Sample/$entry
      -- CP-element group 201: 	 branch_block_stmt_1327/call_stmt_1562_to_assign_stmt_1573/call_stmt_1562_Sample/crr
      -- CP-element group 201: 	 branch_block_stmt_1327/call_stmt_1562_to_assign_stmt_1573/call_stmt_1562_Update/$entry
      -- CP-element group 201: 	 branch_block_stmt_1327/call_stmt_1562_to_assign_stmt_1573/call_stmt_1562_Update/ccr
      -- 
    phi_stmt_1553_ack_3595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1553_ack_0, ack => maxPool3D_CP_2619_elements(201)); -- 
    crr_3069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(201), ack => call_stmt_1562_call_req_0); -- 
    ccr_3074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(201), ack => call_stmt_1562_call_req_1); -- 
    -- CP-element group 202:  merge  transition  place  output  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	54 
    -- CP-element group 202: 	59 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	61 
    -- CP-element group 202:  members (14) 
      -- CP-element group 202: 	 branch_block_stmt_1327/assign_stmt_1599_to_assign_stmt_1603__entry__
      -- CP-element group 202: 	 branch_block_stmt_1327/assign_stmt_1589_to_assign_stmt_1594__exit__
      -- CP-element group 202: 	 branch_block_stmt_1327/assign_stmt_1589_to_assign_stmt_1594__entry__
      -- CP-element group 202: 	 branch_block_stmt_1327/merge_stmt_1582__exit__
      -- CP-element group 202: 	 branch_block_stmt_1327/assign_stmt_1589_to_assign_stmt_1594/$entry
      -- CP-element group 202: 	 branch_block_stmt_1327/assign_stmt_1589_to_assign_stmt_1594/$exit
      -- CP-element group 202: 	 branch_block_stmt_1327/assign_stmt_1599_to_assign_stmt_1603/$entry
      -- CP-element group 202: 	 branch_block_stmt_1327/assign_stmt_1599_to_assign_stmt_1603/WPIPE_maxpool_output_pipe_1596_sample_start_
      -- CP-element group 202: 	 branch_block_stmt_1327/assign_stmt_1599_to_assign_stmt_1603/WPIPE_maxpool_output_pipe_1596_Sample/$entry
      -- CP-element group 202: 	 branch_block_stmt_1327/assign_stmt_1599_to_assign_stmt_1603/WPIPE_maxpool_output_pipe_1596_Sample/req
      -- CP-element group 202: 	 branch_block_stmt_1327/merge_stmt_1582_PhiReqMerge
      -- CP-element group 202: 	 branch_block_stmt_1327/merge_stmt_1582_PhiAck/$entry
      -- CP-element group 202: 	 branch_block_stmt_1327/merge_stmt_1582_PhiAck/$exit
      -- CP-element group 202: 	 branch_block_stmt_1327/merge_stmt_1582_PhiAck/dummy
      -- 
    req_3108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2619_elements(202), ack => WPIPE_maxpool_output_pipe_1596_inst_req_0); -- 
    maxPool3D_CP_2619_elements(202) <= OrReduce(maxPool3D_CP_2619_elements(54) & maxPool3D_CP_2619_elements(59));
    maxPool3D_do_while_stmt_1646_terminator_3447: loop_terminator -- 
      generic map (name => " maxPool3D_do_while_stmt_1646_terminator_3447", max_iterations_in_flight =>15) 
      port map(loop_body_exit => maxPool3D_CP_2619_elements(76),loop_continue => maxPool3D_CP_2619_elements(181),loop_terminate => maxPool3D_CP_2619_elements(180),loop_back => maxPool3D_CP_2619_elements(74),loop_exit => maxPool3D_CP_2619_elements(73),clk => clk, reset => reset); -- 
    phi_stmt_1648_phi_seq_3237_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= maxPool3D_CP_2619_elements(89);
      maxPool3D_CP_2619_elements(94)<= src_sample_reqs(0);
      src_sample_acks(0)  <= maxPool3D_CP_2619_elements(98);
      maxPool3D_CP_2619_elements(95)<= src_update_reqs(0);
      src_update_acks(0)  <= maxPool3D_CP_2619_elements(99);
      maxPool3D_CP_2619_elements(90) <= phi_mux_reqs(0);
      triggers(1)  <= maxPool3D_CP_2619_elements(91);
      maxPool3D_CP_2619_elements(100)<= src_sample_reqs(1);
      src_sample_acks(1)  <= maxPool3D_CP_2619_elements(100);
      maxPool3D_CP_2619_elements(101)<= src_update_reqs(1);
      src_update_acks(1)  <= maxPool3D_CP_2619_elements(102);
      maxPool3D_CP_2619_elements(92) <= phi_mux_reqs(1);
      phi_stmt_1648_phi_seq_3237 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1648_phi_seq_3237") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => maxPool3D_CP_2619_elements(81), 
          phi_sample_ack => maxPool3D_CP_2619_elements(87), 
          phi_update_req => maxPool3D_CP_2619_elements(83), 
          phi_update_ack => maxPool3D_CP_2619_elements(88), 
          phi_mux_ack => maxPool3D_CP_2619_elements(93), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1653_phi_seq_3281_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= maxPool3D_CP_2619_elements(110);
      maxPool3D_CP_2619_elements(115)<= src_sample_reqs(0);
      src_sample_acks(0)  <= maxPool3D_CP_2619_elements(119);
      maxPool3D_CP_2619_elements(116)<= src_update_reqs(0);
      src_update_acks(0)  <= maxPool3D_CP_2619_elements(120);
      maxPool3D_CP_2619_elements(111) <= phi_mux_reqs(0);
      triggers(1)  <= maxPool3D_CP_2619_elements(112);
      maxPool3D_CP_2619_elements(121)<= src_sample_reqs(1);
      src_sample_acks(1)  <= maxPool3D_CP_2619_elements(121);
      maxPool3D_CP_2619_elements(122)<= src_update_reqs(1);
      src_update_acks(1)  <= maxPool3D_CP_2619_elements(123);
      maxPool3D_CP_2619_elements(113) <= phi_mux_reqs(1);
      phi_stmt_1653_phi_seq_3281 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1653_phi_seq_3281") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => maxPool3D_CP_2619_elements(106), 
          phi_sample_ack => maxPool3D_CP_2619_elements(107), 
          phi_update_req => maxPool3D_CP_2619_elements(108), 
          phi_update_ack => maxPool3D_CP_2619_elements(109), 
          phi_mux_ack => maxPool3D_CP_2619_elements(114), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1658_phi_seq_3325_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= maxPool3D_CP_2619_elements(131);
      maxPool3D_CP_2619_elements(136)<= src_sample_reqs(0);
      src_sample_acks(0)  <= maxPool3D_CP_2619_elements(140);
      maxPool3D_CP_2619_elements(137)<= src_update_reqs(0);
      src_update_acks(0)  <= maxPool3D_CP_2619_elements(141);
      maxPool3D_CP_2619_elements(132) <= phi_mux_reqs(0);
      triggers(1)  <= maxPool3D_CP_2619_elements(133);
      maxPool3D_CP_2619_elements(142)<= src_sample_reqs(1);
      src_sample_acks(1)  <= maxPool3D_CP_2619_elements(142);
      maxPool3D_CP_2619_elements(143)<= src_update_reqs(1);
      src_update_acks(1)  <= maxPool3D_CP_2619_elements(144);
      maxPool3D_CP_2619_elements(134) <= phi_mux_reqs(1);
      phi_stmt_1658_phi_seq_3325 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1658_phi_seq_3325") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => maxPool3D_CP_2619_elements(127), 
          phi_sample_ack => maxPool3D_CP_2619_elements(128), 
          phi_update_req => maxPool3D_CP_2619_elements(129), 
          phi_update_ack => maxPool3D_CP_2619_elements(130), 
          phi_mux_ack => maxPool3D_CP_2619_elements(135), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_3189_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= maxPool3D_CP_2619_elements(77);
        preds(1)  <= maxPool3D_CP_2619_elements(78);
        entry_tmerge_3189 : transition_merge -- 
          generic map(name => " entry_tmerge_3189")
          port map (preds => preds, symbol_out => maxPool3D_CP_2619_elements(79));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal NOT_u1_u1_1808_wire : std_logic_vector(0 downto 0);
    signal add114_1685 : std_logic_vector(31 downto 0);
    signal add116_1695 : std_logic_vector(31 downto 0);
    signal add129_1711 : std_logic_vector(31 downto 0);
    signal add132_1721 : std_logic_vector(31 downto 0);
    signal add139_1726 : std_logic_vector(31 downto 0);
    signal add13_1377 : std_logic_vector(15 downto 0);
    signal add143_1731 : std_logic_vector(31 downto 0);
    signal add146_1736 : std_logic_vector(31 downto 0);
    signal add23_1402 : std_logic_vector(15 downto 0);
    signal add33_1427 : std_logic_vector(15 downto 0);
    signal add43_1452 : std_logic_vector(31 downto 0);
    signal add53_1477 : std_logic_vector(15 downto 0);
    signal add98_1627 : std_logic_vector(31 downto 0);
    signal add_1352 : std_logic_vector(31 downto 0);
    signal call11_1368 : std_logic_vector(7 downto 0);
    signal call147_1743 : std_logic_vector(7 downto 0);
    signal call16_1380 : std_logic_vector(7 downto 0);
    signal call21_1393 : std_logic_vector(7 downto 0);
    signal call26_1405 : std_logic_vector(7 downto 0);
    signal call2_1343 : std_logic_vector(7 downto 0);
    signal call31_1418 : std_logic_vector(7 downto 0);
    signal call36_1430 : std_logic_vector(7 downto 0);
    signal call41_1443 : std_logic_vector(7 downto 0);
    signal call46_1455 : std_logic_vector(7 downto 0);
    signal call51_1468 : std_logic_vector(7 downto 0);
    signal call6_1355 : std_logic_vector(7 downto 0);
    signal call_1330 : std_logic_vector(7 downto 0);
    signal chlx_x0_1658 : std_logic_vector(15 downto 0);
    signal chlx_x0_at_entry_1640 : std_logic_vector(15 downto 0);
    signal chlx_x1_1773 : std_logic_vector(15 downto 0);
    signal cmp154_1754 : std_logic_vector(0 downto 0);
    signal cmp162_1778 : std_logic_vector(0 downto 0);
    signal cmp172_1802 : std_logic_vector(0 downto 0);
    signal cmp186_1498 : std_logic_vector(0 downto 0);
    signal colx_x1_1653 : std_logic_vector(15 downto 0);
    signal colx_x1_1749_delayed_1_0_1761 : std_logic_vector(15 downto 0);
    signal colx_x1_at_entry_1635 : std_logic_vector(15 downto 0);
    signal colx_x2_1797 : std_logic_vector(15 downto 0);
    signal conv104_1667 : std_logic_vector(31 downto 0);
    signal conv108_1671 : std_logic_vector(31 downto 0);
    signal conv110_1616 : std_logic_vector(31 downto 0);
    signal conv112_1675 : std_logic_vector(31 downto 0);
    signal conv12_1372 : std_logic_vector(15 downto 0);
    signal conv179_1827 : std_logic_vector(31 downto 0);
    signal conv182_1831 : std_logic_vector(31 downto 0);
    signal conv19_1384 : std_logic_vector(15 downto 0);
    signal conv1_1334 : std_logic_vector(31 downto 0);
    signal conv22_1397 : std_logic_vector(15 downto 0);
    signal conv29_1409 : std_logic_vector(15 downto 0);
    signal conv32_1422 : std_logic_vector(15 downto 0);
    signal conv39_1434 : std_logic_vector(31 downto 0);
    signal conv3_1347 : std_logic_vector(31 downto 0);
    signal conv42_1447 : std_logic_vector(31 downto 0);
    signal conv49_1459 : std_logic_vector(15 downto 0);
    signal conv52_1472 : std_logic_vector(15 downto 0);
    signal conv59_1482 : std_logic_vector(31 downto 0);
    signal conv95_1608 : std_logic_vector(31 downto 0);
    signal conv97_1612 : std_logic_vector(31 downto 0);
    signal conv9_1359 : std_logic_vector(15 downto 0);
    signal exitcond1_1573 : std_logic_vector(0 downto 0);
    signal iNsTr_14_1537 : std_logic_vector(63 downto 0);
    signal iNsTr_24_1553 : std_logic_vector(63 downto 0);
    signal inc149_1749 : std_logic_vector(15 downto 0);
    signal inc157_1758 : std_logic_vector(15 downto 0);
    signal inc157x_xcolx_x1_1766 : std_logic_vector(15 downto 0);
    signal inc166_1782 : std_logic_vector(15 downto 0);
    signal inc166x_xrowx_x1_1790 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_1568 : std_logic_vector(63 downto 0);
    signal mul113_1680 : std_logic_vector(31 downto 0);
    signal mul115_1690 : std_logic_vector(31 downto 0);
    signal mul128_1706 : std_logic_vector(31 downto 0);
    signal mul130_1622 : std_logic_vector(31 downto 0);
    signal mul180_1836 : std_logic_vector(31 downto 0);
    signal mul183_1841 : std_logic_vector(31 downto 0);
    signal mul62_1492 : std_logic_vector(31 downto 0);
    signal mul86_1594 : std_logic_vector(15 downto 0);
    signal mul_1487 : std_logic_vector(31 downto 0);
    signal rowx_x1_1648 : std_logic_vector(15 downto 0);
    signal rowx_x1_1770_delayed_2_0_1785 : std_logic_vector(15 downto 0);
    signal rowx_x1_at_entry_1630 : std_logic_vector(15 downto 0);
    signal shl10_1365 : std_logic_vector(15 downto 0);
    signal shl117_1701 : std_logic_vector(31 downto 0);
    signal shl131_1716 : std_logic_vector(31 downto 0);
    signal shl20_1390 : std_logic_vector(15 downto 0);
    signal shl30_1415 : std_logic_vector(15 downto 0);
    signal shl40_1440 : std_logic_vector(31 downto 0);
    signal shl50_1465 : std_logic_vector(15 downto 0);
    signal shl_1340 : std_logic_vector(31 downto 0);
    signal shr79184_1589 : std_logic_vector(15 downto 0);
    signal tmp189_1515 : std_logic_vector(31 downto 0);
    signal tmp190_1521 : std_logic_vector(31 downto 0);
    signal tmp190x_xop_1533 : std_logic_vector(31 downto 0);
    signal tmp191_1527 : std_logic_vector(0 downto 0);
    signal tmp194_1550 : std_logic_vector(63 downto 0);
    signal tmp_1510 : std_logic_vector(31 downto 0);
    signal type_cast_1338_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1363_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1388_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1413_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1438_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1463_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1496_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1519_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1525_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1531_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1541_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1548_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1557_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1559_wire : std_logic_vector(63 downto 0);
    signal type_cast_1566_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1587_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1598_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1602_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1620_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1651_wire : std_logic_vector(15 downto 0);
    signal type_cast_1656_wire : std_logic_vector(15 downto 0);
    signal type_cast_1661_wire : std_logic_vector(15 downto 0);
    signal type_cast_1699_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1747_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1770_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1794_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1817_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1821_wire_constant : std_logic_vector(7 downto 0);
    signal whilex_xbody_whilex_xend_taken_1805 : std_logic_vector(0 downto 0);
    signal xx_xop_1543 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    chlx_x0_at_entry_1640 <= "0000000000000000";
    colx_x1_at_entry_1635 <= "0000000000000000";
    rowx_x1_at_entry_1630 <= "0000000000000000";
    type_cast_1338_wire_constant <= "00000000000000000000000000001000";
    type_cast_1363_wire_constant <= "0000000000001000";
    type_cast_1388_wire_constant <= "0000000000001000";
    type_cast_1413_wire_constant <= "0000000000001000";
    type_cast_1438_wire_constant <= "00000000000000000000000000001000";
    type_cast_1463_wire_constant <= "0000000000001000";
    type_cast_1496_wire_constant <= "00000000000000000000000000001111";
    type_cast_1519_wire_constant <= "00000000000000000000000000000100";
    type_cast_1525_wire_constant <= "00000000000000000000000000000001";
    type_cast_1531_wire_constant <= "11111111111111111111111111111111";
    type_cast_1541_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1548_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1557_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1566_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1587_wire_constant <= "0000000000000100";
    type_cast_1598_wire_constant <= "11111111";
    type_cast_1602_wire_constant <= "11111111";
    type_cast_1620_wire_constant <= "00000000000000000000000000000001";
    type_cast_1699_wire_constant <= "00000000000000000000000000000010";
    type_cast_1747_wire_constant <= "0000000000000001";
    type_cast_1770_wire_constant <= "0000000000000000";
    type_cast_1794_wire_constant <= "0000000000000000";
    type_cast_1817_wire_constant <= "11111111";
    type_cast_1821_wire_constant <= "11111111";
    phi_stmt_1553: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1557_wire_constant & type_cast_1559_wire;
      req <= phi_stmt_1553_req_0 & phi_stmt_1553_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1553",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1553_ack_0,
          idata => idata,
          odata => iNsTr_24_1553,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1553
    phi_stmt_1648: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1651_wire & rowx_x1_at_entry_1630;
      req <= phi_stmt_1648_req_0 & phi_stmt_1648_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1648",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1648_ack_0,
          idata => idata,
          odata => rowx_x1_1648,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1648
    phi_stmt_1653: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1656_wire & colx_x1_at_entry_1635;
      req <= phi_stmt_1653_req_0 & phi_stmt_1653_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1653",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1653_ack_0,
          idata => idata,
          odata => colx_x1_1653,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1653
    phi_stmt_1658: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1661_wire & chlx_x0_at_entry_1640;
      req <= phi_stmt_1658_req_0 & phi_stmt_1658_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1658",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1658_ack_0,
          idata => idata,
          odata => chlx_x0_1658,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1658
    -- flow-through select operator MUX_1549_inst
    tmp194_1550 <= xx_xop_1543 when (tmp191_1527(0) /=  '0') else type_cast_1548_wire_constant;
    -- flow-through select operator MUX_1772_inst
    chlx_x1_1773 <= type_cast_1770_wire_constant when (cmp154_1754(0) /=  '0') else inc149_1749;
    -- flow-through select operator MUX_1796_inst
    colx_x2_1797 <= type_cast_1794_wire_constant when (cmp162_1778(0) /=  '0') else inc157x_xcolx_x1_1766;
    W_colx_x1_1749_delayed_1_0_1759_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_colx_x1_1749_delayed_1_0_1759_inst_req_0;
      W_colx_x1_1749_delayed_1_0_1759_inst_ack_0<= wack(0);
      rreq(0) <= W_colx_x1_1749_delayed_1_0_1759_inst_req_1;
      W_colx_x1_1749_delayed_1_0_1759_inst_ack_1<= rack(0);
      W_colx_x1_1749_delayed_1_0_1759_inst : InterlockBuffer generic map ( -- 
        name => "W_colx_x1_1749_delayed_1_0_1759_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => colx_x1_1653,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => colx_x1_1749_delayed_1_0_1761,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rowx_x1_1770_delayed_2_0_1783_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rowx_x1_1770_delayed_2_0_1783_inst_req_0;
      W_rowx_x1_1770_delayed_2_0_1783_inst_ack_0<= wack(0);
      rreq(0) <= W_rowx_x1_1770_delayed_2_0_1783_inst_req_1;
      W_rowx_x1_1770_delayed_2_0_1783_inst_ack_1<= rack(0);
      W_rowx_x1_1770_delayed_2_0_1783_inst : InterlockBuffer generic map ( -- 
        name => "W_rowx_x1_1770_delayed_2_0_1783_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rowx_x1_1648,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rowx_x1_1770_delayed_2_0_1785,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_whilex_xbody_whilex_xend_taken_1803_inst
    process(cmp172_1802) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := cmp172_1802(0 downto 0);
      whilex_xbody_whilex_xend_taken_1805 <= tmp_var; -- 
    end process;
    type_cast_1333_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1333_inst_req_0;
      type_cast_1333_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1333_inst_req_1;
      type_cast_1333_inst_ack_1<= rack(0);
      type_cast_1333_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1333_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1330,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1_1334,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1346_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1346_inst_req_0;
      type_cast_1346_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1346_inst_req_1;
      type_cast_1346_inst_ack_1<= rack(0);
      type_cast_1346_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1346_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_1343,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_1347,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1358_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1358_inst_req_0;
      type_cast_1358_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1358_inst_req_1;
      type_cast_1358_inst_ack_1<= rack(0);
      type_cast_1358_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1358_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call6_1355,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv9_1359,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1371_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1371_inst_req_0;
      type_cast_1371_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1371_inst_req_1;
      type_cast_1371_inst_ack_1<= rack(0);
      type_cast_1371_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1371_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call11_1368,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv12_1372,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1383_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1383_inst_req_0;
      type_cast_1383_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1383_inst_req_1;
      type_cast_1383_inst_ack_1<= rack(0);
      type_cast_1383_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1383_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_1380,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv19_1384,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1396_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1396_inst_req_0;
      type_cast_1396_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1396_inst_req_1;
      type_cast_1396_inst_ack_1<= rack(0);
      type_cast_1396_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1396_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call21_1393,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv22_1397,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1408_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1408_inst_req_0;
      type_cast_1408_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1408_inst_req_1;
      type_cast_1408_inst_ack_1<= rack(0);
      type_cast_1408_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1408_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call26_1405,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_1409,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1421_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1421_inst_req_0;
      type_cast_1421_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1421_inst_req_1;
      type_cast_1421_inst_ack_1<= rack(0);
      type_cast_1421_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1421_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call31_1418,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv32_1422,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1433_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1433_inst_req_0;
      type_cast_1433_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1433_inst_req_1;
      type_cast_1433_inst_ack_1<= rack(0);
      type_cast_1433_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1433_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call36_1430,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv39_1434,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1446_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1446_inst_req_0;
      type_cast_1446_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1446_inst_req_1;
      type_cast_1446_inst_ack_1<= rack(0);
      type_cast_1446_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1446_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_1443,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv42_1447,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1458_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1458_inst_req_0;
      type_cast_1458_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1458_inst_req_1;
      type_cast_1458_inst_ack_1<= rack(0);
      type_cast_1458_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1458_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_1455,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv49_1459,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1471_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1471_inst_req_0;
      type_cast_1471_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1471_inst_req_1;
      type_cast_1471_inst_ack_1<= rack(0);
      type_cast_1471_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1471_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call51_1468,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv52_1472,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1481_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1481_inst_req_0;
      type_cast_1481_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1481_inst_req_1;
      type_cast_1481_inst_ack_1<= rack(0);
      type_cast_1481_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1481_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_1402,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv59_1482,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1536_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1536_inst_req_0;
      type_cast_1536_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1536_inst_req_1;
      type_cast_1536_inst_ack_1<= rack(0);
      type_cast_1536_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1536_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp190x_xop_1533,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_14_1537,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1559_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1559_inst_req_0;
      type_cast_1559_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1559_inst_req_1;
      type_cast_1559_inst_ack_1<= rack(0);
      type_cast_1559_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1559_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1568,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1559_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1607_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1607_inst_req_0;
      type_cast_1607_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1607_inst_req_1;
      type_cast_1607_inst_ack_1<= rack(0);
      type_cast_1607_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1607_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr79184_1589,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_1608,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1611_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1611_inst_req_0;
      type_cast_1611_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1611_inst_req_1;
      type_cast_1611_inst_ack_1<= rack(0);
      type_cast_1611_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1611_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul86_1594,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv97_1612,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1615_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1615_inst_req_0;
      type_cast_1615_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1615_inst_req_1;
      type_cast_1615_inst_ack_1<= rack(0);
      type_cast_1615_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1615_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add33_1427,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv110_1616,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1651_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1651_inst_req_0;
      type_cast_1651_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1651_inst_req_1;
      type_cast_1651_inst_ack_1<= rack(0);
      type_cast_1651_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1651_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc166x_xrowx_x1_1790,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1651_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1656_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1656_inst_req_0;
      type_cast_1656_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1656_inst_req_1;
      type_cast_1656_inst_ack_1<= rack(0);
      type_cast_1656_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1656_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => colx_x2_1797,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1656_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1661_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1661_inst_req_0;
      type_cast_1661_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1661_inst_req_1;
      type_cast_1661_inst_ack_1<= rack(0);
      type_cast_1661_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1661_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => chlx_x1_1773,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1661_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1666_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1666_inst_req_0;
      type_cast_1666_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1666_inst_req_1;
      type_cast_1666_inst_ack_1<= rack(0);
      type_cast_1666_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1666_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => chlx_x0_1658,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv104_1667,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1670_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1670_inst_req_0;
      type_cast_1670_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1670_inst_req_1;
      type_cast_1670_inst_ack_1<= rack(0);
      type_cast_1670_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1670_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => colx_x1_1653,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv108_1671,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1674_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1674_inst_req_0;
      type_cast_1674_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1674_inst_req_1;
      type_cast_1674_inst_ack_1<= rack(0);
      type_cast_1674_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1674_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rowx_x1_1648,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv112_1675,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1757_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1757_inst_req_0;
      type_cast_1757_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1757_inst_req_1;
      type_cast_1757_inst_ack_1<= rack(0);
      type_cast_1757_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1757_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp154_1754,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc157_1758,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1781_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1781_inst_req_0;
      type_cast_1781_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1781_inst_req_1;
      type_cast_1781_inst_ack_1<= rack(0);
      type_cast_1781_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1781_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp162_1778,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc166_1782,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1826_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1826_inst_req_0;
      type_cast_1826_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1826_inst_req_1;
      type_cast_1826_inst_ack_1<= rack(0);
      type_cast_1826_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1826_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add13_1377,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv179_1827,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1830_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1830_inst_req_0;
      type_cast_1830_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1830_inst_req_1;
      type_cast_1830_inst_ack_1<= rack(0);
      type_cast_1830_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1830_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add53_1477,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv182_1831,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_1646_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_1808_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1646_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1646_branch_req_0,
          ack0 => do_while_stmt_1646_branch_ack_0,
          ack1 => do_while_stmt_1646_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1499_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp186_1498;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1499_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1499_branch_req_0,
          ack0 => if_stmt_1499_branch_ack_0,
          ack1 => if_stmt_1499_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1574_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_1573;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1574_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1574_branch_req_0,
          ack0 => if_stmt_1574_branch_ack_0,
          ack1 => if_stmt_1574_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1809_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= whilex_xbody_whilex_xend_taken_1805;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1809_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1809_branch_req_0,
          ack0 => if_stmt_1809_branch_ack_0,
          ack1 => if_stmt_1809_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1748_inst
    process(chlx_x0_1658) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(chlx_x0_1658, type_cast_1747_wire_constant, tmp_var);
      inc149_1749 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1765_inst
    process(inc157_1758, colx_x1_1749_delayed_1_0_1761) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc157_1758, colx_x1_1749_delayed_1_0_1761, tmp_var);
      inc157x_xcolx_x1_1766 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1789_inst
    process(inc166_1782, rowx_x1_1770_delayed_2_0_1785) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc166_1782, rowx_x1_1770_delayed_2_0_1785, tmp_var);
      inc166x_xrowx_x1_1790 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1532_inst
    process(tmp190_1521) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp190_1521, type_cast_1531_wire_constant, tmp_var);
      tmp190x_xop_1533 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1626_inst
    process(conv97_1612, conv95_1608) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv97_1612, conv95_1608, tmp_var);
      add98_1627 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1684_inst
    process(conv108_1671, mul113_1680) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv108_1671, mul113_1680, tmp_var);
      add114_1685 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1694_inst
    process(mul115_1690, conv104_1667) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul115_1690, conv104_1667, tmp_var);
      add116_1695 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1710_inst
    process(conv108_1671, mul128_1706) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv108_1671, mul128_1706, tmp_var);
      add129_1711 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1720_inst
    process(shl131_1716, conv104_1667) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl131_1716, conv104_1667, tmp_var);
      add132_1721 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1725_inst
    process(add132_1721, conv95_1608) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add132_1721, conv95_1608, tmp_var);
      add139_1726 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1730_inst
    process(add132_1721, conv97_1612) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add132_1721, conv97_1612, tmp_var);
      add143_1731 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1735_inst
    process(add98_1627, add132_1721) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add98_1627, add132_1721, tmp_var);
      add146_1736 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1542_inst
    process(iNsTr_14_1537) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_14_1537, type_cast_1541_wire_constant, tmp_var);
      xx_xop_1543 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1567_inst
    process(iNsTr_24_1553) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_24_1553, type_cast_1566_wire_constant, tmp_var);
      indvarx_xnext_1568 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1753_inst
    process(inc149_1749, shr79184_1589) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc149_1749, shr79184_1589, tmp_var);
      cmp154_1754 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1777_inst
    process(inc157x_xcolx_x1_1766, add33_1427) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc157x_xcolx_x1_1766, add33_1427, tmp_var);
      cmp162_1778 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1801_inst
    process(inc166x_xrowx_x1_1790, add13_1377) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc166x_xrowx_x1_1790, add13_1377, tmp_var);
      cmp172_1802 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1572_inst
    process(indvarx_xnext_1568, tmp194_1550) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1568, tmp194_1550, tmp_var);
      exitcond1_1573 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_1588_inst
    process(add53_1477) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add53_1477, type_cast_1587_wire_constant, tmp_var);
      shr79184_1589 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1520_inst
    process(tmp189_1515) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp189_1515, type_cast_1519_wire_constant, tmp_var);
      tmp190_1521 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1593_inst
    process(shr79184_1589, add23_1402) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(shr79184_1589, add23_1402, tmp_var);
      mul86_1594 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1486_inst
    process(conv59_1482, add_1352) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv59_1482, add_1352, tmp_var);
      mul_1487 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1491_inst
    process(mul_1487, add43_1452) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_1487, add43_1452, tmp_var);
      mul62_1492 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1509_inst
    process(add_1352, add43_1452) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_1352, add43_1452, tmp_var);
      tmp_1510 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1514_inst
    process(tmp_1510, conv59_1482) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp_1510, conv59_1482, tmp_var);
      tmp189_1515 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1679_inst
    process(conv112_1675, conv110_1616) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv112_1675, conv110_1616, tmp_var);
      mul113_1680 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1689_inst
    process(add114_1685, conv95_1608) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add114_1685, conv95_1608, tmp_var);
      mul115_1690 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1705_inst
    process(conv112_1675, conv59_1482) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv112_1675, conv59_1482, tmp_var);
      mul128_1706 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1715_inst
    process(mul130_1622, add129_1711) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul130_1622, add129_1711, tmp_var);
      shl131_1716 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1835_inst
    process(conv110_1616, conv179_1827) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv110_1616, conv179_1827, tmp_var);
      mul180_1836 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1840_inst
    process(mul180_1836, conv182_1831) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul180_1836, conv182_1831, tmp_var);
      mul183_1841 <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1808_inst
    process(cmp172_1802) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp172_1802, tmp_var);
      NOT_u1_u1_1808_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u16_u16_1376_inst
    process(shl10_1365, conv12_1372) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl10_1365, conv12_1372, tmp_var);
      add13_1377 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1401_inst
    process(shl20_1390, conv22_1397) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl20_1390, conv22_1397, tmp_var);
      add23_1402 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1426_inst
    process(shl30_1415, conv32_1422) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl30_1415, conv32_1422, tmp_var);
      add33_1427 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1476_inst
    process(shl50_1465, conv52_1472) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl50_1465, conv52_1472, tmp_var);
      add53_1477 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1351_inst
    process(shl_1340, conv3_1347) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_1340, conv3_1347, tmp_var);
      add_1352 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1451_inst
    process(shl40_1440, conv42_1447) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl40_1440, conv42_1447, tmp_var);
      add43_1452 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_1364_inst
    process(conv9_1359) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv9_1359, type_cast_1363_wire_constant, tmp_var);
      shl10_1365 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_1389_inst
    process(conv19_1384) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv19_1384, type_cast_1388_wire_constant, tmp_var);
      shl20_1390 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_1414_inst
    process(conv29_1409) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv29_1409, type_cast_1413_wire_constant, tmp_var);
      shl30_1415 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_1464_inst
    process(conv49_1459) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv49_1459, type_cast_1463_wire_constant, tmp_var);
      shl50_1465 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1339_inst
    process(conv1_1334) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1_1334, type_cast_1338_wire_constant, tmp_var);
      shl_1340 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1439_inst
    process(conv39_1434) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv39_1434, type_cast_1438_wire_constant, tmp_var);
      shl40_1440 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1621_inst
    process(conv95_1608) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv95_1608, type_cast_1620_wire_constant, tmp_var);
      mul130_1622 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1700_inst
    process(add116_1695) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add116_1695, type_cast_1699_wire_constant, tmp_var);
      shl117_1701 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1497_inst
    process(mul62_1492) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul62_1492, type_cast_1496_wire_constant, tmp_var);
      cmp186_1498 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1526_inst
    process(tmp190_1521) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp190_1521, type_cast_1525_wire_constant, tmp_var);
      tmp191_1527 <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_maxpool_input_pipe_1329_inst RPIPE_maxpool_input_pipe_1342_inst RPIPE_maxpool_input_pipe_1354_inst RPIPE_maxpool_input_pipe_1367_inst RPIPE_maxpool_input_pipe_1379_inst RPIPE_maxpool_input_pipe_1392_inst RPIPE_maxpool_input_pipe_1404_inst RPIPE_maxpool_input_pipe_1417_inst RPIPE_maxpool_input_pipe_1429_inst RPIPE_maxpool_input_pipe_1442_inst RPIPE_maxpool_input_pipe_1454_inst RPIPE_maxpool_input_pipe_1467_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(95 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 11 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 11 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 11 downto 0);
      signal guard_vector : std_logic_vector( 11 downto 0);
      constant outBUFs : IntegerArray(11 downto 0) := (11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(11 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false);
      constant guardBuffering: IntegerArray(11 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2);
      -- 
    begin -- 
      reqL_unguarded(11) <= RPIPE_maxpool_input_pipe_1329_inst_req_0;
      reqL_unguarded(10) <= RPIPE_maxpool_input_pipe_1342_inst_req_0;
      reqL_unguarded(9) <= RPIPE_maxpool_input_pipe_1354_inst_req_0;
      reqL_unguarded(8) <= RPIPE_maxpool_input_pipe_1367_inst_req_0;
      reqL_unguarded(7) <= RPIPE_maxpool_input_pipe_1379_inst_req_0;
      reqL_unguarded(6) <= RPIPE_maxpool_input_pipe_1392_inst_req_0;
      reqL_unguarded(5) <= RPIPE_maxpool_input_pipe_1404_inst_req_0;
      reqL_unguarded(4) <= RPIPE_maxpool_input_pipe_1417_inst_req_0;
      reqL_unguarded(3) <= RPIPE_maxpool_input_pipe_1429_inst_req_0;
      reqL_unguarded(2) <= RPIPE_maxpool_input_pipe_1442_inst_req_0;
      reqL_unguarded(1) <= RPIPE_maxpool_input_pipe_1454_inst_req_0;
      reqL_unguarded(0) <= RPIPE_maxpool_input_pipe_1467_inst_req_0;
      RPIPE_maxpool_input_pipe_1329_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_maxpool_input_pipe_1342_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_maxpool_input_pipe_1354_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_maxpool_input_pipe_1367_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_maxpool_input_pipe_1379_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_maxpool_input_pipe_1392_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_maxpool_input_pipe_1404_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_maxpool_input_pipe_1417_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_maxpool_input_pipe_1429_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_maxpool_input_pipe_1442_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_maxpool_input_pipe_1454_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_maxpool_input_pipe_1467_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(11) <= RPIPE_maxpool_input_pipe_1329_inst_req_1;
      reqR_unguarded(10) <= RPIPE_maxpool_input_pipe_1342_inst_req_1;
      reqR_unguarded(9) <= RPIPE_maxpool_input_pipe_1354_inst_req_1;
      reqR_unguarded(8) <= RPIPE_maxpool_input_pipe_1367_inst_req_1;
      reqR_unguarded(7) <= RPIPE_maxpool_input_pipe_1379_inst_req_1;
      reqR_unguarded(6) <= RPIPE_maxpool_input_pipe_1392_inst_req_1;
      reqR_unguarded(5) <= RPIPE_maxpool_input_pipe_1404_inst_req_1;
      reqR_unguarded(4) <= RPIPE_maxpool_input_pipe_1417_inst_req_1;
      reqR_unguarded(3) <= RPIPE_maxpool_input_pipe_1429_inst_req_1;
      reqR_unguarded(2) <= RPIPE_maxpool_input_pipe_1442_inst_req_1;
      reqR_unguarded(1) <= RPIPE_maxpool_input_pipe_1454_inst_req_1;
      reqR_unguarded(0) <= RPIPE_maxpool_input_pipe_1467_inst_req_1;
      RPIPE_maxpool_input_pipe_1329_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_maxpool_input_pipe_1342_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_maxpool_input_pipe_1354_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_maxpool_input_pipe_1367_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_maxpool_input_pipe_1379_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_maxpool_input_pipe_1392_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_maxpool_input_pipe_1404_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_maxpool_input_pipe_1417_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_maxpool_input_pipe_1429_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_maxpool_input_pipe_1442_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_maxpool_input_pipe_1454_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_maxpool_input_pipe_1467_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      call_1330 <= data_out(95 downto 88);
      call2_1343 <= data_out(87 downto 80);
      call6_1355 <= data_out(79 downto 72);
      call11_1368 <= data_out(71 downto 64);
      call16_1380 <= data_out(63 downto 56);
      call21_1393 <= data_out(55 downto 48);
      call26_1405 <= data_out(47 downto 40);
      call31_1418 <= data_out(39 downto 32);
      call36_1430 <= data_out(31 downto 24);
      call41_1443 <= data_out(23 downto 16);
      call46_1455 <= data_out(15 downto 8);
      call51_1468 <= data_out(7 downto 0);
      maxpool_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "maxpool_input_pipe_read_0_gI", nreqs => 12, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      maxpool_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "maxpool_input_pipe_read_0", data_width => 8,  num_reqs => 12,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => maxpool_input_pipe_pipe_read_req(0),
          oack => maxpool_input_pipe_pipe_read_ack(0),
          odata => maxpool_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_maxpool_output_pipe_1815_inst WPIPE_maxpool_output_pipe_1819_inst WPIPE_maxpool_output_pipe_1600_inst WPIPE_maxpool_output_pipe_1596_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 3 downto 0);
      signal update_req, update_ack : BooleanArray( 3 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 3 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      sample_req_unguarded(3) <= WPIPE_maxpool_output_pipe_1815_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_maxpool_output_pipe_1819_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1600_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1596_inst_req_0;
      WPIPE_maxpool_output_pipe_1815_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_1819_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_1600_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1596_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(3) <= WPIPE_maxpool_output_pipe_1815_inst_req_1;
      update_req_unguarded(2) <= WPIPE_maxpool_output_pipe_1819_inst_req_1;
      update_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1600_inst_req_1;
      update_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1596_inst_req_1;
      WPIPE_maxpool_output_pipe_1815_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_1819_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_1600_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1596_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      data_in <= type_cast_1817_wire_constant & type_cast_1821_wire_constant & type_cast_1602_wire_constant & type_cast_1598_wire_constant;
      maxpool_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "maxpool_output_pipe_write_0_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      maxpool_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "maxpool_output_pipe", data_width => 8, num_reqs => 4, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => maxpool_output_pipe_pipe_write_req(0),
          oack => maxpool_output_pipe_pipe_write_ack(0),
          odata => maxpool_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_1562_call 
    fill_T_call_group_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1562_call_req_0;
      call_stmt_1562_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1562_call_req_1;
      call_stmt_1562_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      fill_T_call_group_0_gI: SplitGuardInterface generic map(name => "fill_T_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= iNsTr_24_1553;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 64,
        owidth => 64,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => fill_T_call_reqs(0),
          ackR => fill_T_call_acks(0),
          dataR => fill_T_call_data(63 downto 0),
          tagR => fill_T_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => fill_T_return_acks(0), -- cross-over
          ackL => fill_T_return_reqs(0), -- cross-over
          tagL => fill_T_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1743_call 
    maxPool4_call_group_1: Block -- 
      signal data_in: std_logic_vector(159 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 17);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1743_call_req_0;
      call_stmt_1743_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1743_call_req_1;
      call_stmt_1743_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      maxPool4_call_group_1_gI: SplitGuardInterface generic map(name => "maxPool4_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= shl117_1701 & add132_1721 & add139_1726 & add143_1731 & add146_1736;
      call147_1743 <= data_out(7 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 160,
        owidth => 160,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => maxPool4_call_reqs(0),
          ackR => maxPool4_call_acks(0),
          dataR => maxPool4_call_data(159 downto 0),
          tagR => maxPool4_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 8,
          owidth => 8,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => maxPool4_return_acks(0), -- cross-over
          ackL => maxPool4_return_reqs(0), -- cross-over
          dataL => maxPool4_return_data(7 downto 0),
          tagL => maxPool4_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_1843_call 
    sendB_call_group_2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1843_call_req_0;
      call_stmt_1843_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1843_call_req_1;
      call_stmt_1843_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      sendB_call_group_2_gI: SplitGuardInterface generic map(name => "sendB_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= mul183_1841;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 32,
        owidth => 32,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => sendB_call_reqs(0),
          ackR => sendB_call_acks(0),
          dataR => sendB_call_data(31 downto 0),
          tagR => sendB_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => sendB_return_acks(0), -- cross-over
          ackL => sendB_return_reqs(0), -- cross-over
          tagL => sendB_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- 
  end Block; -- data_path
  -- 
end maxPool3D_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity maxPool4 is -- 
  generic (tag_length : integer); 
  port ( -- 
    addr : in  std_logic_vector(31 downto 0);
    addr1 : in  std_logic_vector(31 downto 0);
    addr2 : in  std_logic_vector(31 downto 0);
    addr3 : in  std_logic_vector(31 downto 0);
    addr4 : in  std_logic_vector(31 downto 0);
    output : out  std_logic_vector(7 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(255 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity maxPool4;
architecture maxPool4_arch of maxPool4 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 160)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 8)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal addr_buffer :  std_logic_vector(31 downto 0);
  signal addr_update_enable: Boolean;
  signal addr1_buffer :  std_logic_vector(31 downto 0);
  signal addr1_update_enable: Boolean;
  signal addr2_buffer :  std_logic_vector(31 downto 0);
  signal addr2_update_enable: Boolean;
  signal addr3_buffer :  std_logic_vector(31 downto 0);
  signal addr3_update_enable: Boolean;
  signal addr4_buffer :  std_logic_vector(31 downto 0);
  signal addr4_update_enable: Boolean;
  -- output port buffer signals
  signal output_buffer :  std_logic_vector(7 downto 0);
  signal output_update_enable: Boolean;
  signal maxPool4_CP_307_start: Boolean;
  signal maxPool4_CP_307_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal slice_222_inst_ack_1 : boolean;
  signal CONCAT_u32_u64_1047_inst_ack_1 : boolean;
  signal slice_222_inst_req_1 : boolean;
  signal slice_210_inst_ack_1 : boolean;
  signal slice_234_inst_ack_0 : boolean;
  signal slice_374_inst_req_0 : boolean;
  signal slice_242_inst_req_1 : boolean;
  signal slice_242_inst_req_0 : boolean;
  signal slice_238_inst_ack_1 : boolean;
  signal slice_238_inst_req_1 : boolean;
  signal slice_210_inst_req_1 : boolean;
  signal slice_270_inst_req_1 : boolean;
  signal slice_246_inst_ack_0 : boolean;
  signal slice_234_inst_req_0 : boolean;
  signal slice_246_inst_req_0 : boolean;
  signal slice_214_inst_ack_1 : boolean;
  signal slice_222_inst_ack_0 : boolean;
  signal ptr_deref_1036_store_0_req_1 : boolean;
  signal slice_214_inst_req_1 : boolean;
  signal slice_382_inst_req_1 : boolean;
  signal ptr_deref_1036_store_0_ack_0 : boolean;
  signal slice_226_inst_ack_0 : boolean;
  signal slice_238_inst_ack_0 : boolean;
  signal slice_226_inst_req_0 : boolean;
  signal ptr_deref_1036_store_0_ack_1 : boolean;
  signal ptr_deref_1036_store_0_req_0 : boolean;
  signal slice_238_inst_req_0 : boolean;
  signal slice_222_inst_req_0 : boolean;
  signal slice_374_inst_ack_0 : boolean;
  signal addr_of_1030_final_reg_req_1 : boolean;
  signal slice_214_inst_ack_0 : boolean;
  signal slice_234_inst_ack_1 : boolean;
  signal slice_218_inst_req_1 : boolean;
  signal slice_234_inst_req_1 : boolean;
  signal slice_250_inst_ack_0 : boolean;
  signal CONCAT_u32_u64_1073_inst_req_1 : boolean;
  signal slice_254_inst_ack_1 : boolean;
  signal slice_250_inst_ack_1 : boolean;
  signal slice_250_inst_req_1 : boolean;
  signal slice_258_inst_ack_1 : boolean;
  signal slice_254_inst_req_1 : boolean;
  signal slice_214_inst_req_0 : boolean;
  signal slice_374_inst_req_1 : boolean;
  signal slice_250_inst_req_0 : boolean;
  signal slice_270_inst_ack_1 : boolean;
  signal slice_374_inst_ack_1 : boolean;
  signal slice_274_inst_ack_0 : boolean;
  signal ptr_deref_1062_store_0_req_0 : boolean;
  signal addr_of_1030_final_reg_ack_1 : boolean;
  signal slice_262_inst_req_1 : boolean;
  signal addr_of_1030_final_reg_req_0 : boolean;
  signal slice_266_inst_ack_1 : boolean;
  signal addr_of_1030_final_reg_ack_0 : boolean;
  signal slice_270_inst_ack_0 : boolean;
  signal slice_262_inst_ack_0 : boolean;
  signal slice_270_inst_req_0 : boolean;
  signal ptr_deref_1062_store_0_ack_0 : boolean;
  signal slice_218_inst_ack_1 : boolean;
  signal slice_266_inst_req_1 : boolean;
  signal slice_382_inst_ack_1 : boolean;
  signal slice_262_inst_ack_1 : boolean;
  signal CONCAT_u32_u64_1073_inst_ack_1 : boolean;
  signal slice_262_inst_req_0 : boolean;
  signal slice_274_inst_req_0 : boolean;
  signal slice_258_inst_req_1 : boolean;
  signal slice_254_inst_ack_0 : boolean;
  signal W_myptr6_1055_delayed_8_0_1058_inst_req_1 : boolean;
  signal ptr_deref_117_load_0_req_0 : boolean;
  signal ptr_deref_117_load_0_ack_0 : boolean;
  signal ptr_deref_117_load_0_req_1 : boolean;
  signal ptr_deref_117_load_0_ack_1 : boolean;
  signal slice_254_inst_req_0 : boolean;
  signal slice_210_inst_ack_0 : boolean;
  signal slice_242_inst_ack_0 : boolean;
  signal slice_210_inst_req_0 : boolean;
  signal slice_218_inst_ack_0 : boolean;
  signal slice_230_inst_ack_1 : boolean;
  signal slice_230_inst_req_1 : boolean;
  signal slice_266_inst_ack_0 : boolean;
  signal slice_266_inst_req_0 : boolean;
  signal slice_246_inst_ack_1 : boolean;
  signal slice_230_inst_ack_0 : boolean;
  signal slice_230_inst_req_0 : boolean;
  signal slice_258_inst_ack_0 : boolean;
  signal slice_258_inst_req_0 : boolean;
  signal slice_226_inst_ack_1 : boolean;
  signal slice_226_inst_req_1 : boolean;
  signal array_obj_ref_87_index_offset_req_0 : boolean;
  signal array_obj_ref_87_index_offset_ack_0 : boolean;
  signal slice_218_inst_req_0 : boolean;
  signal array_obj_ref_87_index_offset_req_1 : boolean;
  signal array_obj_ref_87_index_offset_ack_1 : boolean;
  signal slice_242_inst_ack_1 : boolean;
  signal slice_246_inst_req_1 : boolean;
  signal addr_of_88_final_reg_req_0 : boolean;
  signal addr_of_88_final_reg_ack_0 : boolean;
  signal addr_of_88_final_reg_req_1 : boolean;
  signal addr_of_88_final_reg_ack_1 : boolean;
  signal array_obj_ref_94_index_offset_req_0 : boolean;
  signal array_obj_ref_94_index_offset_ack_0 : boolean;
  signal array_obj_ref_94_index_offset_req_1 : boolean;
  signal array_obj_ref_94_index_offset_ack_1 : boolean;
  signal addr_of_95_final_reg_req_0 : boolean;
  signal addr_of_95_final_reg_ack_0 : boolean;
  signal addr_of_95_final_reg_req_1 : boolean;
  signal addr_of_95_final_reg_ack_1 : boolean;
  signal W_myptr5_1032_delayed_8_0_1032_inst_req_0 : boolean;
  signal W_myptr5_1032_delayed_8_0_1032_inst_ack_0 : boolean;
  signal array_obj_ref_101_index_offset_req_0 : boolean;
  signal array_obj_ref_101_index_offset_ack_0 : boolean;
  signal array_obj_ref_101_index_offset_req_1 : boolean;
  signal array_obj_ref_101_index_offset_ack_1 : boolean;
  signal addr_of_102_final_reg_req_0 : boolean;
  signal addr_of_102_final_reg_ack_0 : boolean;
  signal addr_of_102_final_reg_req_1 : boolean;
  signal addr_of_102_final_reg_ack_1 : boolean;
  signal W_myptr5_1032_delayed_8_0_1032_inst_req_1 : boolean;
  signal array_obj_ref_108_index_offset_req_0 : boolean;
  signal array_obj_ref_108_index_offset_ack_0 : boolean;
  signal W_myptr5_1032_delayed_8_0_1032_inst_ack_1 : boolean;
  signal array_obj_ref_108_index_offset_req_1 : boolean;
  signal array_obj_ref_108_index_offset_ack_1 : boolean;
  signal addr_of_109_final_reg_req_0 : boolean;
  signal addr_of_109_final_reg_ack_0 : boolean;
  signal W_myptr6_1055_delayed_8_0_1058_inst_req_0 : boolean;
  signal addr_of_109_final_reg_req_1 : boolean;
  signal addr_of_109_final_reg_ack_1 : boolean;
  signal slice_378_inst_req_0 : boolean;
  signal slice_378_inst_ack_0 : boolean;
  signal ptr_deref_113_load_0_req_0 : boolean;
  signal ptr_deref_113_load_0_ack_0 : boolean;
  signal ptr_deref_113_load_0_req_1 : boolean;
  signal ptr_deref_113_load_0_ack_1 : boolean;
  signal slice_378_inst_req_1 : boolean;
  signal W_myptr6_1055_delayed_8_0_1058_inst_ack_0 : boolean;
  signal array_obj_ref_1055_index_offset_req_0 : boolean;
  signal CONCAT_u32_u64_1047_inst_req_0 : boolean;
  signal array_obj_ref_1055_index_offset_ack_0 : boolean;
  signal ptr_deref_121_load_0_req_0 : boolean;
  signal ptr_deref_121_load_0_ack_0 : boolean;
  signal ptr_deref_121_load_0_req_1 : boolean;
  signal ptr_deref_121_load_0_ack_1 : boolean;
  signal slice_378_inst_ack_1 : boolean;
  signal addr_of_1082_final_reg_ack_0 : boolean;
  signal array_obj_ref_1055_index_offset_req_1 : boolean;
  signal slice_274_inst_req_1 : boolean;
  signal slice_274_inst_ack_1 : boolean;
  signal CONCAT_u32_u64_1047_inst_ack_0 : boolean;
  signal ptr_deref_125_load_0_req_0 : boolean;
  signal array_obj_ref_1055_index_offset_ack_1 : boolean;
  signal ptr_deref_125_load_0_ack_0 : boolean;
  signal ptr_deref_125_load_0_req_1 : boolean;
  signal ptr_deref_125_load_0_ack_1 : boolean;
  signal CONCAT_u32_u64_1047_inst_req_1 : boolean;
  signal slice_130_inst_req_0 : boolean;
  signal slice_130_inst_ack_0 : boolean;
  signal slice_130_inst_req_1 : boolean;
  signal slice_130_inst_ack_1 : boolean;
  signal slice_134_inst_req_0 : boolean;
  signal slice_134_inst_ack_0 : boolean;
  signal slice_134_inst_req_1 : boolean;
  signal slice_134_inst_ack_1 : boolean;
  signal slice_138_inst_req_0 : boolean;
  signal slice_138_inst_ack_0 : boolean;
  signal slice_382_inst_req_0 : boolean;
  signal slice_138_inst_req_1 : boolean;
  signal slice_138_inst_ack_1 : boolean;
  signal slice_382_inst_ack_0 : boolean;
  signal slice_142_inst_req_0 : boolean;
  signal slice_142_inst_ack_0 : boolean;
  signal slice_142_inst_req_1 : boolean;
  signal slice_142_inst_ack_1 : boolean;
  signal slice_146_inst_req_0 : boolean;
  signal slice_146_inst_ack_0 : boolean;
  signal slice_146_inst_req_1 : boolean;
  signal slice_146_inst_ack_1 : boolean;
  signal slice_150_inst_req_0 : boolean;
  signal slice_150_inst_ack_0 : boolean;
  signal slice_150_inst_req_1 : boolean;
  signal slice_150_inst_ack_1 : boolean;
  signal slice_154_inst_req_0 : boolean;
  signal slice_154_inst_ack_0 : boolean;
  signal slice_154_inst_req_1 : boolean;
  signal slice_154_inst_ack_1 : boolean;
  signal slice_158_inst_req_0 : boolean;
  signal slice_158_inst_ack_0 : boolean;
  signal slice_158_inst_req_1 : boolean;
  signal slice_158_inst_ack_1 : boolean;
  signal slice_162_inst_req_0 : boolean;
  signal slice_162_inst_ack_0 : boolean;
  signal slice_162_inst_req_1 : boolean;
  signal slice_162_inst_ack_1 : boolean;
  signal slice_166_inst_req_0 : boolean;
  signal slice_166_inst_ack_0 : boolean;
  signal slice_166_inst_req_1 : boolean;
  signal slice_166_inst_ack_1 : boolean;
  signal slice_170_inst_req_0 : boolean;
  signal slice_170_inst_ack_0 : boolean;
  signal slice_170_inst_req_1 : boolean;
  signal slice_170_inst_ack_1 : boolean;
  signal slice_174_inst_req_0 : boolean;
  signal slice_174_inst_ack_0 : boolean;
  signal slice_174_inst_req_1 : boolean;
  signal slice_174_inst_ack_1 : boolean;
  signal slice_178_inst_req_0 : boolean;
  signal slice_178_inst_ack_0 : boolean;
  signal slice_178_inst_req_1 : boolean;
  signal slice_178_inst_ack_1 : boolean;
  signal slice_182_inst_req_0 : boolean;
  signal slice_182_inst_ack_0 : boolean;
  signal slice_182_inst_req_1 : boolean;
  signal slice_182_inst_ack_1 : boolean;
  signal slice_186_inst_req_0 : boolean;
  signal slice_186_inst_ack_0 : boolean;
  signal slice_186_inst_req_1 : boolean;
  signal slice_186_inst_ack_1 : boolean;
  signal slice_190_inst_req_0 : boolean;
  signal slice_190_inst_ack_0 : boolean;
  signal slice_190_inst_req_1 : boolean;
  signal slice_190_inst_ack_1 : boolean;
  signal slice_194_inst_req_0 : boolean;
  signal slice_194_inst_ack_0 : boolean;
  signal slice_194_inst_req_1 : boolean;
  signal slice_194_inst_ack_1 : boolean;
  signal slice_198_inst_req_0 : boolean;
  signal slice_198_inst_ack_0 : boolean;
  signal slice_198_inst_req_1 : boolean;
  signal slice_198_inst_ack_1 : boolean;
  signal slice_202_inst_req_0 : boolean;
  signal slice_202_inst_ack_0 : boolean;
  signal slice_202_inst_req_1 : boolean;
  signal slice_202_inst_ack_1 : boolean;
  signal slice_206_inst_req_0 : boolean;
  signal slice_206_inst_ack_0 : boolean;
  signal slice_206_inst_req_1 : boolean;
  signal slice_206_inst_ack_1 : boolean;
  signal addr_of_1082_final_reg_req_1 : boolean;
  signal addr_of_1082_final_reg_ack_1 : boolean;
  signal slice_370_inst_ack_1 : boolean;
  signal slice_278_inst_req_0 : boolean;
  signal slice_278_inst_ack_0 : boolean;
  signal addr_of_1056_final_reg_ack_1 : boolean;
  signal slice_278_inst_req_1 : boolean;
  signal slice_278_inst_ack_1 : boolean;
  signal array_obj_ref_1081_index_offset_ack_1 : boolean;
  signal slice_370_inst_req_1 : boolean;
  signal slice_282_inst_req_0 : boolean;
  signal slice_282_inst_ack_0 : boolean;
  signal addr_of_1056_final_reg_req_1 : boolean;
  signal slice_282_inst_req_1 : boolean;
  signal slice_282_inst_ack_1 : boolean;
  signal array_obj_ref_1081_index_offset_req_1 : boolean;
  signal ptr_deref_1062_store_0_ack_1 : boolean;
  signal slice_286_inst_req_0 : boolean;
  signal slice_286_inst_ack_0 : boolean;
  signal slice_286_inst_req_1 : boolean;
  signal slice_286_inst_ack_1 : boolean;
  signal array_obj_ref_1029_index_offset_ack_1 : boolean;
  signal slice_290_inst_req_0 : boolean;
  signal slice_290_inst_ack_0 : boolean;
  signal slice_290_inst_req_1 : boolean;
  signal slice_290_inst_ack_1 : boolean;
  signal array_obj_ref_1029_index_offset_req_1 : boolean;
  signal ptr_deref_1062_store_0_req_1 : boolean;
  signal slice_370_inst_ack_0 : boolean;
  signal slice_294_inst_req_0 : boolean;
  signal slice_294_inst_ack_0 : boolean;
  signal addr_of_1056_final_reg_ack_0 : boolean;
  signal slice_294_inst_req_1 : boolean;
  signal slice_294_inst_ack_1 : boolean;
  signal array_obj_ref_1081_index_offset_ack_0 : boolean;
  signal slice_370_inst_req_0 : boolean;
  signal array_obj_ref_1029_index_offset_ack_0 : boolean;
  signal slice_298_inst_req_0 : boolean;
  signal slice_298_inst_ack_0 : boolean;
  signal addr_of_1056_final_reg_req_0 : boolean;
  signal slice_298_inst_req_1 : boolean;
  signal slice_298_inst_ack_1 : boolean;
  signal array_obj_ref_1081_index_offset_req_0 : boolean;
  signal array_obj_ref_1029_index_offset_req_0 : boolean;
  signal slice_302_inst_req_0 : boolean;
  signal slice_302_inst_ack_0 : boolean;
  signal slice_302_inst_req_1 : boolean;
  signal slice_302_inst_ack_1 : boolean;
  signal addr_of_1082_final_reg_req_0 : boolean;
  signal slice_306_inst_req_0 : boolean;
  signal slice_306_inst_ack_0 : boolean;
  signal slice_306_inst_req_1 : boolean;
  signal slice_306_inst_ack_1 : boolean;
  signal slice_310_inst_req_0 : boolean;
  signal slice_310_inst_ack_0 : boolean;
  signal slice_310_inst_req_1 : boolean;
  signal slice_310_inst_ack_1 : boolean;
  signal CONCAT_u32_u64_1073_inst_ack_0 : boolean;
  signal slice_366_inst_ack_1 : boolean;
  signal slice_314_inst_req_0 : boolean;
  signal slice_314_inst_ack_0 : boolean;
  signal slice_366_inst_req_1 : boolean;
  signal slice_314_inst_req_1 : boolean;
  signal slice_314_inst_ack_1 : boolean;
  signal slice_318_inst_req_0 : boolean;
  signal slice_318_inst_ack_0 : boolean;
  signal slice_366_inst_ack_0 : boolean;
  signal slice_318_inst_req_1 : boolean;
  signal slice_318_inst_ack_1 : boolean;
  signal CONCAT_u32_u64_1073_inst_req_0 : boolean;
  signal slice_366_inst_req_0 : boolean;
  signal W_myptr6_1055_delayed_8_0_1058_inst_ack_1 : boolean;
  signal slice_322_inst_req_0 : boolean;
  signal slice_322_inst_ack_0 : boolean;
  signal slice_322_inst_req_1 : boolean;
  signal slice_322_inst_ack_1 : boolean;
  signal slice_326_inst_req_0 : boolean;
  signal slice_326_inst_ack_0 : boolean;
  signal slice_326_inst_req_1 : boolean;
  signal slice_326_inst_ack_1 : boolean;
  signal slice_330_inst_req_0 : boolean;
  signal slice_330_inst_ack_0 : boolean;
  signal slice_330_inst_req_1 : boolean;
  signal slice_330_inst_ack_1 : boolean;
  signal slice_334_inst_req_0 : boolean;
  signal slice_334_inst_ack_0 : boolean;
  signal slice_334_inst_req_1 : boolean;
  signal slice_334_inst_ack_1 : boolean;
  signal slice_338_inst_req_0 : boolean;
  signal slice_338_inst_ack_0 : boolean;
  signal slice_338_inst_req_1 : boolean;
  signal slice_338_inst_ack_1 : boolean;
  signal slice_342_inst_req_0 : boolean;
  signal slice_342_inst_ack_0 : boolean;
  signal slice_342_inst_req_1 : boolean;
  signal slice_342_inst_ack_1 : boolean;
  signal slice_346_inst_req_0 : boolean;
  signal slice_346_inst_ack_0 : boolean;
  signal slice_346_inst_req_1 : boolean;
  signal slice_346_inst_ack_1 : boolean;
  signal slice_350_inst_req_0 : boolean;
  signal slice_350_inst_ack_0 : boolean;
  signal slice_350_inst_req_1 : boolean;
  signal slice_350_inst_ack_1 : boolean;
  signal slice_354_inst_req_0 : boolean;
  signal slice_354_inst_ack_0 : boolean;
  signal slice_354_inst_req_1 : boolean;
  signal slice_354_inst_ack_1 : boolean;
  signal slice_358_inst_req_0 : boolean;
  signal slice_358_inst_ack_0 : boolean;
  signal slice_358_inst_req_1 : boolean;
  signal slice_358_inst_ack_1 : boolean;
  signal slice_362_inst_req_0 : boolean;
  signal slice_362_inst_ack_0 : boolean;
  signal slice_362_inst_req_1 : boolean;
  signal slice_362_inst_ack_1 : boolean;
  signal W_myptr7_1078_delayed_8_0_1084_inst_req_0 : boolean;
  signal W_myptr7_1078_delayed_8_0_1084_inst_ack_0 : boolean;
  signal W_myptr7_1078_delayed_8_0_1084_inst_req_1 : boolean;
  signal W_myptr7_1078_delayed_8_0_1084_inst_ack_1 : boolean;
  signal CONCAT_u32_u64_1099_inst_req_0 : boolean;
  signal CONCAT_u32_u64_1099_inst_ack_0 : boolean;
  signal CONCAT_u32_u64_1099_inst_req_1 : boolean;
  signal CONCAT_u32_u64_1099_inst_ack_1 : boolean;
  signal ptr_deref_1088_store_0_req_0 : boolean;
  signal ptr_deref_1088_store_0_ack_0 : boolean;
  signal ptr_deref_1088_store_0_req_1 : boolean;
  signal ptr_deref_1088_store_0_ack_1 : boolean;
  signal array_obj_ref_1107_index_offset_req_0 : boolean;
  signal array_obj_ref_1107_index_offset_ack_0 : boolean;
  signal array_obj_ref_1107_index_offset_req_1 : boolean;
  signal array_obj_ref_1107_index_offset_ack_1 : boolean;
  signal addr_of_1108_final_reg_req_0 : boolean;
  signal addr_of_1108_final_reg_ack_0 : boolean;
  signal addr_of_1108_final_reg_req_1 : boolean;
  signal addr_of_1108_final_reg_ack_1 : boolean;
  signal W_myptr8_1101_delayed_8_0_1110_inst_req_0 : boolean;
  signal W_myptr8_1101_delayed_8_0_1110_inst_ack_0 : boolean;
  signal W_myptr8_1101_delayed_8_0_1110_inst_req_1 : boolean;
  signal W_myptr8_1101_delayed_8_0_1110_inst_ack_1 : boolean;
  signal CONCAT_u32_u64_1125_inst_req_0 : boolean;
  signal CONCAT_u32_u64_1125_inst_ack_0 : boolean;
  signal CONCAT_u32_u64_1125_inst_req_1 : boolean;
  signal CONCAT_u32_u64_1125_inst_ack_1 : boolean;
  signal ptr_deref_1114_store_0_req_0 : boolean;
  signal ptr_deref_1114_store_0_ack_0 : boolean;
  signal ptr_deref_1114_store_0_req_1 : boolean;
  signal ptr_deref_1114_store_0_ack_1 : boolean;
  signal type_cast_1129_inst_req_0 : boolean;
  signal type_cast_1129_inst_ack_0 : boolean;
  signal type_cast_1129_inst_req_1 : boolean;
  signal type_cast_1129_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "maxPool4_input_buffer", -- 
      buffer_size => 2,
      bypass_flag => false,
      data_width => tag_length + 160) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= addr;
  addr_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(63 downto 32) <= addr1;
  addr1_buffer <= in_buffer_data_out(63 downto 32);
  in_buffer_data_in(95 downto 64) <= addr2;
  addr2_buffer <= in_buffer_data_out(95 downto 64);
  in_buffer_data_in(127 downto 96) <= addr3;
  addr3_buffer <= in_buffer_data_out(127 downto 96);
  in_buffer_data_in(159 downto 128) <= addr4;
  addr4_buffer <= in_buffer_data_out(159 downto 128);
  in_buffer_data_in(tag_length + 159 downto 160) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 159 downto 160);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 1,6 => 15);
    constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1,6 => 15);
    constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 7); -- 
  begin -- 
    preds <= addr_update_enable & addr1_update_enable & addr2_update_enable & addr3_update_enable & addr4_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  maxPool4_CP_307_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "maxPool4_out_buffer", -- 
      buffer_size => 2,
      full_rate => false,
      data_width => tag_length + 8) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(7 downto 0) <= output_buffer;
  output <= out_buffer_data_out(7 downto 0);
  out_buffer_data_in(tag_length + 7 downto 8) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 7 downto 8);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 15);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= maxPool4_CP_307_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  output_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 25) := "output_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_output_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => output_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 15,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= maxPool4_CP_307_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= maxPool4_CP_307_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  maxPool4_CP_307: Block -- control-path 
    signal maxPool4_CP_307_elements: BooleanArray(398 downto 0);
    -- 
  begin -- 
    maxPool4_CP_307_elements(0) <= maxPool4_CP_307_start;
    maxPool4_CP_307_symbol <= maxPool4_CP_307_elements(398);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	9 
    -- CP-element group 1: 	10 
    -- CP-element group 1: 	11 
    -- CP-element group 1: 	16 
    -- CP-element group 1: 	17 
    -- CP-element group 1: 	18 
    -- CP-element group 1: 	23 
    -- CP-element group 1: 	24 
    -- CP-element group 1: 	25 
    -- CP-element group 1: 	30 
    -- CP-element group 1: 	31 
    -- CP-element group 1: 	32 
    -- CP-element group 1: 	309 
    -- CP-element group 1: 	310 
    -- CP-element group 1: 	311 
    -- CP-element group 1: 	328 
    -- CP-element group 1: 	329 
    -- CP-element group 1: 	330 
    -- CP-element group 1: 	347 
    -- CP-element group 1: 	348 
    -- CP-element group 1: 	349 
    -- CP-element group 1: 	366 
    -- CP-element group 1: 	367 
    -- CP-element group 1: 	368 
    -- CP-element group 1:  members (105) 
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1081_index_scale_1/$entry
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1029_index_scaled_1
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1081_index_resize_1/index_resize_req
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1081_index_resize_1/$entry
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1081_final_index_sum_regn_Sample/$entry
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1055_final_index_sum_regn_Sample/$entry
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1081_index_scale_1/$exit
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/$entry
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_87_index_resized_1
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_87_index_scaled_1
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_87_index_computed_1
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_87_index_resize_1/$entry
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_87_index_resize_1/$exit
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_87_index_resize_1/index_resize_req
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_87_index_resize_1/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_87_index_scale_1/$entry
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_87_index_scale_1/$exit
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_87_index_scale_1/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_87_index_scale_1/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_87_final_index_sum_regn_Sample/$entry
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_87_final_index_sum_regn_Sample/req
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_94_index_resized_1
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_94_index_scaled_1
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_94_index_computed_1
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_94_index_resize_1/$entry
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_94_index_resize_1/$exit
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_94_index_resize_1/index_resize_req
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_94_index_resize_1/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_94_index_scale_1/$entry
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_94_index_scale_1/$exit
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_94_index_scale_1/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_94_index_scale_1/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1055_index_resized_1
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_94_final_index_sum_regn_Sample/$entry
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_94_final_index_sum_regn_Sample/req
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1055_index_scaled_1
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1055_index_computed_1
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1055_index_resize_1/$entry
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_101_index_resized_1
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_101_index_scaled_1
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_101_index_computed_1
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_101_index_resize_1/$entry
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_101_index_resize_1/$exit
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_101_index_resize_1/index_resize_req
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_101_index_resize_1/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_101_index_scale_1/$entry
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_101_index_scale_1/$exit
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_101_index_scale_1/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_101_index_scale_1/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_101_final_index_sum_regn_Sample/$entry
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_101_final_index_sum_regn_Sample/req
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_108_index_resized_1
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_108_index_scaled_1
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_108_index_computed_1
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1055_index_resize_1/$exit
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_108_index_resize_1/$entry
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_108_index_resize_1/$exit
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_108_index_resize_1/index_resize_req
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_108_index_resize_1/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_108_index_scale_1/$entry
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_108_index_scale_1/$exit
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_108_index_scale_1/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_108_index_scale_1/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1055_index_resize_1/index_resize_req
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_108_final_index_sum_regn_Sample/$entry
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_108_final_index_sum_regn_Sample/req
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1081_index_resize_1/$exit
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1055_index_resize_1/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1055_index_scale_1/$entry
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1055_index_scale_1/$exit
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1055_index_scale_1/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1055_index_scale_1/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1055_final_index_sum_regn_Sample/req
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1081_index_resize_1/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1029_index_resized_1
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1081_index_scale_1/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1081_index_scale_1/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1081_index_computed_1
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1081_index_scaled_1
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1081_index_resized_1
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1081_final_index_sum_regn_Sample/req
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1029_final_index_sum_regn_Sample/req
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1029_final_index_sum_regn_Sample/$entry
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1029_index_scale_1/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1029_index_scale_1/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1029_index_scale_1/$exit
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1029_index_scale_1/$entry
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1029_index_resize_1/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1029_index_resize_1/index_resize_req
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1029_index_resize_1/$exit
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1029_index_resize_1/$entry
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1029_index_computed_1
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1107_index_resized_1
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1107_index_scaled_1
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1107_index_computed_1
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1107_index_resize_1/$entry
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1107_index_resize_1/$exit
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1107_index_resize_1/index_resize_req
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1107_index_resize_1/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1107_index_scale_1/$entry
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1107_index_scale_1/$exit
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1107_index_scale_1/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1107_index_scale_1/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1107_final_index_sum_regn_Sample/$entry
      -- CP-element group 1: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1107_final_index_sum_regn_Sample/req
      -- 
    req_349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(1), ack => array_obj_ref_87_index_offset_req_0); -- 
    req_395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(1), ack => array_obj_ref_94_index_offset_req_0); -- 
    req_441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(1), ack => array_obj_ref_101_index_offset_req_0); -- 
    req_487_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_487_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(1), ack => array_obj_ref_108_index_offset_req_0); -- 
    req_1629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(1), ack => array_obj_ref_1029_index_offset_req_0); -- 
    req_1753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(1), ack => array_obj_ref_1055_index_offset_req_0); -- 
    req_1877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(1), ack => array_obj_ref_1081_index_offset_req_0); -- 
    req_2001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(1), ack => array_obj_ref_1107_index_offset_req_0); -- 
    maxPool4_CP_307_elements(1) <= maxPool4_CP_307_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	311 
    -- CP-element group 2: 	330 
    -- CP-element group 2: 	349 
    -- CP-element group 2: 	368 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	392 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 assign_stmt_89_to_assign_stmt_1130/addr_update_enable
      -- CP-element group 2: 	 assign_stmt_89_to_assign_stmt_1130/addr_update_enable_out
      -- 
    maxPool4_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(311) & maxPool4_CP_307_elements(330) & maxPool4_CP_307_elements(349) & maxPool4_CP_307_elements(368);
      gj_maxPool4_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  join  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: marked-predecessors 
    -- CP-element group 3: 	11 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	393 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 assign_stmt_89_to_assign_stmt_1130/addr1_update_enable
      -- CP-element group 3: 	 assign_stmt_89_to_assign_stmt_1130/addr1_update_enable_out
      -- 
    maxPool4_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 1);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_307_elements(11);
      gj_maxPool4_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  join  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: marked-predecessors 
    -- CP-element group 4: 	18 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	394 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 assign_stmt_89_to_assign_stmt_1130/addr2_update_enable
      -- CP-element group 4: 	 assign_stmt_89_to_assign_stmt_1130/addr2_update_enable_out
      -- 
    maxPool4_cp_element_group_4: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 1);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_4"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_307_elements(18);
      gj_maxPool4_cp_element_group_4 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(4), clk => clk, reset => reset); --
    end block;
    -- CP-element group 5:  join  transition  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: marked-predecessors 
    -- CP-element group 5: 	25 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	395 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 assign_stmt_89_to_assign_stmt_1130/addr3_update_enable
      -- CP-element group 5: 	 assign_stmt_89_to_assign_stmt_1130/addr3_update_enable_out
      -- 
    maxPool4_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 1);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_307_elements(25);
      gj_maxPool4_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  join  transition  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	32 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	396 
    -- CP-element group 6:  members (2) 
      -- CP-element group 6: 	 assign_stmt_89_to_assign_stmt_1130/addr4_update_enable
      -- CP-element group 6: 	 assign_stmt_89_to_assign_stmt_1130/addr4_update_enable_out
      -- 
    maxPool4_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 1);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_307_elements(32);
      gj_maxPool4_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	397 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	385 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 assign_stmt_89_to_assign_stmt_1130/output_update_enable
      -- CP-element group 7: 	 assign_stmt_89_to_assign_stmt_1130/output_update_enable_in
      -- 
    maxPool4_CP_307_elements(7) <= maxPool4_CP_307_elements(397);
    -- CP-element group 8:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	12 
    -- CP-element group 8: marked-predecessors 
    -- CP-element group 8: 	13 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	13 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_88_sample_start_
      -- CP-element group 8: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_88_request/$entry
      -- CP-element group 8: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_88_request/req
      -- 
    req_364_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_364_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(8), ack => addr_of_88_final_reg_req_0); -- 
    maxPool4_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(12) & maxPool4_CP_307_elements(13);
      gj_maxPool4_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	1 
    -- CP-element group 9: marked-predecessors 
    -- CP-element group 9: 	14 
    -- CP-element group 9: 	38 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	14 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_88_update_start_
      -- CP-element group 9: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_88_complete/$entry
      -- CP-element group 9: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_88_complete/req
      -- 
    req_369_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_369_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(9), ack => addr_of_88_final_reg_req_1); -- 
    maxPool4_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(1) & maxPool4_CP_307_elements(14) & maxPool4_CP_307_elements(38);
      gj_maxPool4_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	1 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	12 
    -- CP-element group 10: 	13 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_87_final_index_sum_regn_update_start
      -- CP-element group 10: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_87_final_index_sum_regn_Update/$entry
      -- CP-element group 10: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_87_final_index_sum_regn_Update/req
      -- 
    req_354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(10), ack => array_obj_ref_87_index_offset_req_1); -- 
    maxPool4_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(1) & maxPool4_CP_307_elements(12) & maxPool4_CP_307_elements(13);
      gj_maxPool4_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	1 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	391 
    -- CP-element group 11: marked-successors 
    -- CP-element group 11: 	3 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_87_final_index_sum_regn_sample_complete
      -- CP-element group 11: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_87_final_index_sum_regn_Sample/$exit
      -- CP-element group 11: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_87_final_index_sum_regn_Sample/ack
      -- 
    ack_350_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_87_index_offset_ack_0, ack => maxPool4_CP_307_elements(11)); -- 
    -- CP-element group 12:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	8 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	10 
    -- CP-element group 12:  members (8) 
      -- CP-element group 12: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_87_root_address_calculated
      -- CP-element group 12: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_87_offset_calculated
      -- CP-element group 12: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_87_final_index_sum_regn_Update/$exit
      -- CP-element group 12: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_87_final_index_sum_regn_Update/ack
      -- CP-element group 12: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_87_base_plus_offset/$entry
      -- CP-element group 12: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_87_base_plus_offset/$exit
      -- CP-element group 12: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_87_base_plus_offset/sum_rename_req
      -- CP-element group 12: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_87_base_plus_offset/sum_rename_ack
      -- 
    ack_355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_87_index_offset_ack_1, ack => maxPool4_CP_307_elements(12)); -- 
    -- CP-element group 13:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	8 
    -- CP-element group 13: successors 
    -- CP-element group 13: marked-successors 
    -- CP-element group 13: 	8 
    -- CP-element group 13: 	10 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_88_sample_completed_
      -- CP-element group 13: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_88_request/$exit
      -- CP-element group 13: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_88_request/ack
      -- 
    ack_365_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_88_final_reg_ack_0, ack => maxPool4_CP_307_elements(13)); -- 
    -- CP-element group 14:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	9 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	36 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	9 
    -- CP-element group 14:  members (19) 
      -- CP-element group 14: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_88_update_completed_
      -- CP-element group 14: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_88_complete/$exit
      -- CP-element group 14: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_88_complete/ack
      -- CP-element group 14: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_113_base_address_calculated
      -- CP-element group 14: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_113_word_address_calculated
      -- CP-element group 14: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_113_root_address_calculated
      -- CP-element group 14: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_113_base_address_resized
      -- CP-element group 14: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_113_base_addr_resize/$entry
      -- CP-element group 14: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_113_base_addr_resize/$exit
      -- CP-element group 14: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_113_base_addr_resize/base_resize_req
      -- CP-element group 14: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_113_base_addr_resize/base_resize_ack
      -- CP-element group 14: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_113_base_plus_offset/$entry
      -- CP-element group 14: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_113_base_plus_offset/$exit
      -- CP-element group 14: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_113_base_plus_offset/sum_rename_req
      -- CP-element group 14: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_113_base_plus_offset/sum_rename_ack
      -- CP-element group 14: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_113_word_addrgen/$entry
      -- CP-element group 14: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_113_word_addrgen/$exit
      -- CP-element group 14: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_113_word_addrgen/root_register_req
      -- CP-element group 14: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_113_word_addrgen/root_register_ack
      -- 
    ack_370_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_88_final_reg_ack_1, ack => maxPool4_CP_307_elements(14)); -- 
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	19 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	20 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	20 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_95_sample_start_
      -- CP-element group 15: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_95_request/$entry
      -- CP-element group 15: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_95_request/req
      -- 
    req_410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(15), ack => addr_of_95_final_reg_req_0); -- 
    maxPool4_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(19) & maxPool4_CP_307_elements(20);
      gj_maxPool4_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	1 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	21 
    -- CP-element group 16: 	42 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	21 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_95_update_start_
      -- CP-element group 16: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_95_complete/$entry
      -- CP-element group 16: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_95_complete/req
      -- 
    req_415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(16), ack => addr_of_95_final_reg_req_1); -- 
    maxPool4_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(1) & maxPool4_CP_307_elements(21) & maxPool4_CP_307_elements(42);
      gj_maxPool4_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	1 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	19 
    -- CP-element group 17: 	20 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	19 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_94_final_index_sum_regn_update_start
      -- CP-element group 17: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_94_final_index_sum_regn_Update/$entry
      -- CP-element group 17: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_94_final_index_sum_regn_Update/req
      -- 
    req_400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(17), ack => array_obj_ref_94_index_offset_req_1); -- 
    maxPool4_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(1) & maxPool4_CP_307_elements(19) & maxPool4_CP_307_elements(20);
      gj_maxPool4_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	1 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	391 
    -- CP-element group 18: marked-successors 
    -- CP-element group 18: 	4 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_94_final_index_sum_regn_sample_complete
      -- CP-element group 18: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_94_final_index_sum_regn_Sample/$exit
      -- CP-element group 18: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_94_final_index_sum_regn_Sample/ack
      -- 
    ack_396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_94_index_offset_ack_0, ack => maxPool4_CP_307_elements(18)); -- 
    -- CP-element group 19:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	17 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	17 
    -- CP-element group 19:  members (8) 
      -- CP-element group 19: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_94_root_address_calculated
      -- CP-element group 19: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_94_offset_calculated
      -- CP-element group 19: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_94_final_index_sum_regn_Update/$exit
      -- CP-element group 19: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_94_final_index_sum_regn_Update/ack
      -- CP-element group 19: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_94_base_plus_offset/$entry
      -- CP-element group 19: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_94_base_plus_offset/$exit
      -- CP-element group 19: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_94_base_plus_offset/sum_rename_req
      -- CP-element group 19: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_94_base_plus_offset/sum_rename_ack
      -- 
    ack_401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_94_index_offset_ack_1, ack => maxPool4_CP_307_elements(19)); -- 
    -- CP-element group 20:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	15 
    -- CP-element group 20: successors 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	15 
    -- CP-element group 20: 	17 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_95_sample_completed_
      -- CP-element group 20: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_95_request/$exit
      -- CP-element group 20: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_95_request/ack
      -- 
    ack_411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_95_final_reg_ack_0, ack => maxPool4_CP_307_elements(20)); -- 
    -- CP-element group 21:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	16 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	40 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	16 
    -- CP-element group 21:  members (19) 
      -- CP-element group 21: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_117_word_addrgen/root_register_req
      -- CP-element group 21: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_117_word_addrgen/root_register_ack
      -- CP-element group 21: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_95_update_completed_
      -- CP-element group 21: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_95_complete/$exit
      -- CP-element group 21: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_95_complete/ack
      -- CP-element group 21: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_117_base_address_calculated
      -- CP-element group 21: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_117_word_address_calculated
      -- CP-element group 21: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_117_root_address_calculated
      -- CP-element group 21: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_117_base_address_resized
      -- CP-element group 21: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_117_base_addr_resize/$entry
      -- CP-element group 21: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_117_base_addr_resize/$exit
      -- CP-element group 21: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_117_base_addr_resize/base_resize_req
      -- CP-element group 21: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_117_base_addr_resize/base_resize_ack
      -- CP-element group 21: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_117_base_plus_offset/$entry
      -- CP-element group 21: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_117_base_plus_offset/$exit
      -- CP-element group 21: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_117_base_plus_offset/sum_rename_req
      -- CP-element group 21: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_117_base_plus_offset/sum_rename_ack
      -- CP-element group 21: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_117_word_addrgen/$entry
      -- CP-element group 21: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_117_word_addrgen/$exit
      -- 
    ack_416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_95_final_reg_ack_1, ack => maxPool4_CP_307_elements(21)); -- 
    -- CP-element group 22:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	26 
    -- CP-element group 22: marked-predecessors 
    -- CP-element group 22: 	27 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	27 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_102_sample_start_
      -- CP-element group 22: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_102_request/$entry
      -- CP-element group 22: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_102_request/req
      -- 
    req_456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(22), ack => addr_of_102_final_reg_req_0); -- 
    maxPool4_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(26) & maxPool4_CP_307_elements(27);
      gj_maxPool4_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	1 
    -- CP-element group 23: marked-predecessors 
    -- CP-element group 23: 	28 
    -- CP-element group 23: 	46 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	28 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_102_update_start_
      -- CP-element group 23: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_102_complete/$entry
      -- CP-element group 23: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_102_complete/req
      -- 
    req_461_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_461_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(23), ack => addr_of_102_final_reg_req_1); -- 
    maxPool4_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(1) & maxPool4_CP_307_elements(28) & maxPool4_CP_307_elements(46);
      gj_maxPool4_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	1 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	26 
    -- CP-element group 24: 	27 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_101_final_index_sum_regn_update_start
      -- CP-element group 24: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_101_final_index_sum_regn_Update/$entry
      -- CP-element group 24: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_101_final_index_sum_regn_Update/req
      -- 
    req_446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(24), ack => array_obj_ref_101_index_offset_req_1); -- 
    maxPool4_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(1) & maxPool4_CP_307_elements(26) & maxPool4_CP_307_elements(27);
      gj_maxPool4_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	1 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	391 
    -- CP-element group 25: marked-successors 
    -- CP-element group 25: 	5 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_101_final_index_sum_regn_sample_complete
      -- CP-element group 25: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_101_final_index_sum_regn_Sample/$exit
      -- CP-element group 25: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_101_final_index_sum_regn_Sample/ack
      -- 
    ack_442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_101_index_offset_ack_0, ack => maxPool4_CP_307_elements(25)); -- 
    -- CP-element group 26:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	22 
    -- CP-element group 26: marked-successors 
    -- CP-element group 26: 	24 
    -- CP-element group 26:  members (8) 
      -- CP-element group 26: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_101_root_address_calculated
      -- CP-element group 26: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_101_offset_calculated
      -- CP-element group 26: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_101_final_index_sum_regn_Update/$exit
      -- CP-element group 26: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_101_final_index_sum_regn_Update/ack
      -- CP-element group 26: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_101_base_plus_offset/$entry
      -- CP-element group 26: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_101_base_plus_offset/$exit
      -- CP-element group 26: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_101_base_plus_offset/sum_rename_req
      -- CP-element group 26: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_101_base_plus_offset/sum_rename_ack
      -- 
    ack_447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_101_index_offset_ack_1, ack => maxPool4_CP_307_elements(26)); -- 
    -- CP-element group 27:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	22 
    -- CP-element group 27: successors 
    -- CP-element group 27: marked-successors 
    -- CP-element group 27: 	22 
    -- CP-element group 27: 	24 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_102_sample_completed_
      -- CP-element group 27: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_102_request/$exit
      -- CP-element group 27: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_102_request/ack
      -- 
    ack_457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_102_final_reg_ack_0, ack => maxPool4_CP_307_elements(27)); -- 
    -- CP-element group 28:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	23 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	44 
    -- CP-element group 28: marked-successors 
    -- CP-element group 28: 	23 
    -- CP-element group 28:  members (19) 
      -- CP-element group 28: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_102_update_completed_
      -- CP-element group 28: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_102_complete/$exit
      -- CP-element group 28: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_102_complete/ack
      -- CP-element group 28: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_121_base_address_calculated
      -- CP-element group 28: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_121_word_address_calculated
      -- CP-element group 28: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_121_root_address_calculated
      -- CP-element group 28: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_121_base_address_resized
      -- CP-element group 28: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_121_base_addr_resize/$entry
      -- CP-element group 28: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_121_base_addr_resize/$exit
      -- CP-element group 28: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_121_base_addr_resize/base_resize_req
      -- CP-element group 28: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_121_base_addr_resize/base_resize_ack
      -- CP-element group 28: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_121_base_plus_offset/$entry
      -- CP-element group 28: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_121_base_plus_offset/$exit
      -- CP-element group 28: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_121_base_plus_offset/sum_rename_req
      -- CP-element group 28: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_121_base_plus_offset/sum_rename_ack
      -- CP-element group 28: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_121_word_addrgen/$entry
      -- CP-element group 28: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_121_word_addrgen/$exit
      -- CP-element group 28: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_121_word_addrgen/root_register_req
      -- CP-element group 28: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_121_word_addrgen/root_register_ack
      -- 
    ack_462_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_102_final_reg_ack_1, ack => maxPool4_CP_307_elements(28)); -- 
    -- CP-element group 29:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	33 
    -- CP-element group 29: marked-predecessors 
    -- CP-element group 29: 	34 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	34 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_109_sample_start_
      -- CP-element group 29: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_109_request/$entry
      -- CP-element group 29: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_109_request/req
      -- 
    req_502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(29), ack => addr_of_109_final_reg_req_0); -- 
    maxPool4_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(33) & maxPool4_CP_307_elements(34);
      gj_maxPool4_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	1 
    -- CP-element group 30: marked-predecessors 
    -- CP-element group 30: 	35 
    -- CP-element group 30: 	50 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	35 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_109_update_start_
      -- CP-element group 30: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_109_complete/$entry
      -- CP-element group 30: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_109_complete/req
      -- 
    req_507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(30), ack => addr_of_109_final_reg_req_1); -- 
    maxPool4_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(1) & maxPool4_CP_307_elements(35) & maxPool4_CP_307_elements(50);
      gj_maxPool4_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	1 
    -- CP-element group 31: marked-predecessors 
    -- CP-element group 31: 	33 
    -- CP-element group 31: 	34 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_108_final_index_sum_regn_update_start
      -- CP-element group 31: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_108_final_index_sum_regn_Update/$entry
      -- CP-element group 31: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_108_final_index_sum_regn_Update/req
      -- 
    req_492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(31), ack => array_obj_ref_108_index_offset_req_1); -- 
    maxPool4_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(1) & maxPool4_CP_307_elements(33) & maxPool4_CP_307_elements(34);
      gj_maxPool4_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	1 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	391 
    -- CP-element group 32: marked-successors 
    -- CP-element group 32: 	6 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_108_final_index_sum_regn_sample_complete
      -- CP-element group 32: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_108_final_index_sum_regn_Sample/$exit
      -- CP-element group 32: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_108_final_index_sum_regn_Sample/ack
      -- 
    ack_488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_108_index_offset_ack_0, ack => maxPool4_CP_307_elements(32)); -- 
    -- CP-element group 33:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	29 
    -- CP-element group 33: marked-successors 
    -- CP-element group 33: 	31 
    -- CP-element group 33:  members (8) 
      -- CP-element group 33: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_108_root_address_calculated
      -- CP-element group 33: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_108_offset_calculated
      -- CP-element group 33: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_108_final_index_sum_regn_Update/$exit
      -- CP-element group 33: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_108_final_index_sum_regn_Update/ack
      -- CP-element group 33: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_108_base_plus_offset/$entry
      -- CP-element group 33: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_108_base_plus_offset/$exit
      -- CP-element group 33: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_108_base_plus_offset/sum_rename_req
      -- CP-element group 33: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_108_base_plus_offset/sum_rename_ack
      -- 
    ack_493_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_108_index_offset_ack_1, ack => maxPool4_CP_307_elements(33)); -- 
    -- CP-element group 34:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	29 
    -- CP-element group 34: successors 
    -- CP-element group 34: marked-successors 
    -- CP-element group 34: 	29 
    -- CP-element group 34: 	31 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_109_sample_completed_
      -- CP-element group 34: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_109_request/$exit
      -- CP-element group 34: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_109_request/ack
      -- 
    ack_503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_109_final_reg_ack_0, ack => maxPool4_CP_307_elements(34)); -- 
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	30 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	48 
    -- CP-element group 35: marked-successors 
    -- CP-element group 35: 	30 
    -- CP-element group 35:  members (19) 
      -- CP-element group 35: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_125_root_address_calculated
      -- CP-element group 35: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_109_update_completed_
      -- CP-element group 35: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_109_complete/$exit
      -- CP-element group 35: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_109_complete/ack
      -- CP-element group 35: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_125_base_address_calculated
      -- CP-element group 35: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_125_word_address_calculated
      -- CP-element group 35: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_125_base_address_resized
      -- CP-element group 35: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_125_base_addr_resize/$entry
      -- CP-element group 35: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_125_base_addr_resize/$exit
      -- CP-element group 35: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_125_base_addr_resize/base_resize_req
      -- CP-element group 35: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_125_base_addr_resize/base_resize_ack
      -- CP-element group 35: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_125_base_plus_offset/$entry
      -- CP-element group 35: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_125_base_plus_offset/$exit
      -- CP-element group 35: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_125_base_plus_offset/sum_rename_req
      -- CP-element group 35: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_125_base_plus_offset/sum_rename_ack
      -- CP-element group 35: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_125_word_addrgen/$entry
      -- CP-element group 35: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_125_word_addrgen/$exit
      -- CP-element group 35: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_125_word_addrgen/root_register_req
      -- CP-element group 35: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_125_word_addrgen/root_register_ack
      -- 
    ack_508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_109_final_reg_ack_1, ack => maxPool4_CP_307_elements(35)); -- 
    -- CP-element group 36:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	14 
    -- CP-element group 36: marked-predecessors 
    -- CP-element group 36: 	38 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (5) 
      -- CP-element group 36: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_113_sample_start_
      -- CP-element group 36: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_113_Sample/$entry
      -- CP-element group 36: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_113_Sample/word_access_start/$entry
      -- CP-element group 36: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_113_Sample/word_access_start/word_0/$entry
      -- CP-element group 36: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_113_Sample/word_access_start/word_0/rr
      -- 
    rr_541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(36), ack => ptr_deref_113_load_0_req_0); -- 
    maxPool4_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(14) & maxPool4_CP_307_elements(38);
      gj_maxPool4_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	39 
    -- CP-element group 37: 	54 
    -- CP-element group 37: 	58 
    -- CP-element group 37: 	62 
    -- CP-element group 37: 	66 
    -- CP-element group 37: 	70 
    -- CP-element group 37: 	74 
    -- CP-element group 37: 	78 
    -- CP-element group 37: 	82 
    -- CP-element group 37: 	86 
    -- CP-element group 37: 	90 
    -- CP-element group 37: 	94 
    -- CP-element group 37: 	98 
    -- CP-element group 37: 	102 
    -- CP-element group 37: 	106 
    -- CP-element group 37: 	110 
    -- CP-element group 37: 	114 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (5) 
      -- CP-element group 37: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_113_update_start_
      -- CP-element group 37: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_113_Update/$entry
      -- CP-element group 37: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_113_Update/word_access_complete/$entry
      -- CP-element group 37: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_113_Update/word_access_complete/word_0/$entry
      -- CP-element group 37: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_113_Update/word_access_complete/word_0/cr
      -- 
    cr_552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(37), ack => ptr_deref_113_load_0_req_1); -- 
    maxPool4_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(39) & maxPool4_CP_307_elements(54) & maxPool4_CP_307_elements(58) & maxPool4_CP_307_elements(62) & maxPool4_CP_307_elements(66) & maxPool4_CP_307_elements(70) & maxPool4_CP_307_elements(74) & maxPool4_CP_307_elements(78) & maxPool4_CP_307_elements(82) & maxPool4_CP_307_elements(86) & maxPool4_CP_307_elements(90) & maxPool4_CP_307_elements(94) & maxPool4_CP_307_elements(98) & maxPool4_CP_307_elements(102) & maxPool4_CP_307_elements(106) & maxPool4_CP_307_elements(110) & maxPool4_CP_307_elements(114);
      gj_maxPool4_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38: marked-successors 
    -- CP-element group 38: 	9 
    -- CP-element group 38: 	36 
    -- CP-element group 38:  members (5) 
      -- CP-element group 38: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_113_sample_completed_
      -- CP-element group 38: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_113_Sample/$exit
      -- CP-element group 38: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_113_Sample/word_access_start/$exit
      -- CP-element group 38: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_113_Sample/word_access_start/word_0/$exit
      -- CP-element group 38: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_113_Sample/word_access_start/word_0/ra
      -- 
    ra_542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_113_load_0_ack_0, ack => maxPool4_CP_307_elements(38)); -- 
    -- CP-element group 39:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	52 
    -- CP-element group 39: 	56 
    -- CP-element group 39: 	60 
    -- CP-element group 39: 	64 
    -- CP-element group 39: 	68 
    -- CP-element group 39: 	72 
    -- CP-element group 39: 	76 
    -- CP-element group 39: 	80 
    -- CP-element group 39: 	84 
    -- CP-element group 39: 	88 
    -- CP-element group 39: 	92 
    -- CP-element group 39: 	96 
    -- CP-element group 39: 	100 
    -- CP-element group 39: 	104 
    -- CP-element group 39: 	108 
    -- CP-element group 39: 	112 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	37 
    -- CP-element group 39:  members (9) 
      -- CP-element group 39: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_113_update_completed_
      -- CP-element group 39: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_113_Update/$exit
      -- CP-element group 39: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_113_Update/word_access_complete/$exit
      -- CP-element group 39: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_113_Update/word_access_complete/word_0/$exit
      -- CP-element group 39: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_113_Update/word_access_complete/word_0/ca
      -- CP-element group 39: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_113_Update/ptr_deref_113_Merge/$entry
      -- CP-element group 39: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_113_Update/ptr_deref_113_Merge/$exit
      -- CP-element group 39: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_113_Update/ptr_deref_113_Merge/merge_req
      -- CP-element group 39: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_113_Update/ptr_deref_113_Merge/merge_ack
      -- 
    ca_553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_113_load_0_ack_1, ack => maxPool4_CP_307_elements(39)); -- 
    -- CP-element group 40:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	21 
    -- CP-element group 40: marked-predecessors 
    -- CP-element group 40: 	42 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	42 
    -- CP-element group 40:  members (5) 
      -- CP-element group 40: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_117_Sample/$entry
      -- CP-element group 40: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_117_Sample/word_access_start/$entry
      -- CP-element group 40: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_117_Sample/word_access_start/word_0/$entry
      -- CP-element group 40: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_117_Sample/word_access_start/word_0/rr
      -- CP-element group 40: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_117_sample_start_
      -- 
    rr_591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(40), ack => ptr_deref_117_load_0_req_0); -- 
    maxPool4_cp_element_group_40: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_40"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(21) & maxPool4_CP_307_elements(42);
      gj_maxPool4_cp_element_group_40 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(40), clk => clk, reset => reset); --
    end block;
    -- CP-element group 41:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: marked-predecessors 
    -- CP-element group 41: 	43 
    -- CP-element group 41: 	118 
    -- CP-element group 41: 	122 
    -- CP-element group 41: 	126 
    -- CP-element group 41: 	130 
    -- CP-element group 41: 	134 
    -- CP-element group 41: 	138 
    -- CP-element group 41: 	142 
    -- CP-element group 41: 	146 
    -- CP-element group 41: 	150 
    -- CP-element group 41: 	154 
    -- CP-element group 41: 	158 
    -- CP-element group 41: 	162 
    -- CP-element group 41: 	166 
    -- CP-element group 41: 	170 
    -- CP-element group 41: 	174 
    -- CP-element group 41: 	178 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	43 
    -- CP-element group 41:  members (5) 
      -- CP-element group 41: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_117_Update/$entry
      -- CP-element group 41: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_117_Update/word_access_complete/$entry
      -- CP-element group 41: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_117_Update/word_access_complete/word_0/$entry
      -- CP-element group 41: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_117_Update/word_access_complete/word_0/cr
      -- CP-element group 41: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_117_update_start_
      -- 
    cr_602_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_602_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(41), ack => ptr_deref_117_load_0_req_1); -- 
    maxPool4_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(43) & maxPool4_CP_307_elements(118) & maxPool4_CP_307_elements(122) & maxPool4_CP_307_elements(126) & maxPool4_CP_307_elements(130) & maxPool4_CP_307_elements(134) & maxPool4_CP_307_elements(138) & maxPool4_CP_307_elements(142) & maxPool4_CP_307_elements(146) & maxPool4_CP_307_elements(150) & maxPool4_CP_307_elements(154) & maxPool4_CP_307_elements(158) & maxPool4_CP_307_elements(162) & maxPool4_CP_307_elements(166) & maxPool4_CP_307_elements(170) & maxPool4_CP_307_elements(174) & maxPool4_CP_307_elements(178);
      gj_maxPool4_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	40 
    -- CP-element group 42: successors 
    -- CP-element group 42: marked-successors 
    -- CP-element group 42: 	16 
    -- CP-element group 42: 	40 
    -- CP-element group 42:  members (5) 
      -- CP-element group 42: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_117_Sample/$exit
      -- CP-element group 42: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_117_Sample/word_access_start/$exit
      -- CP-element group 42: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_117_Sample/word_access_start/word_0/$exit
      -- CP-element group 42: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_117_Sample/word_access_start/word_0/ra
      -- CP-element group 42: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_117_sample_completed_
      -- 
    ra_592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_117_load_0_ack_0, ack => maxPool4_CP_307_elements(42)); -- 
    -- CP-element group 43:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	41 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	116 
    -- CP-element group 43: 	120 
    -- CP-element group 43: 	124 
    -- CP-element group 43: 	128 
    -- CP-element group 43: 	132 
    -- CP-element group 43: 	136 
    -- CP-element group 43: 	140 
    -- CP-element group 43: 	144 
    -- CP-element group 43: 	148 
    -- CP-element group 43: 	152 
    -- CP-element group 43: 	156 
    -- CP-element group 43: 	160 
    -- CP-element group 43: 	164 
    -- CP-element group 43: 	168 
    -- CP-element group 43: 	172 
    -- CP-element group 43: 	176 
    -- CP-element group 43: marked-successors 
    -- CP-element group 43: 	41 
    -- CP-element group 43:  members (9) 
      -- CP-element group 43: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_117_Update/$exit
      -- CP-element group 43: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_117_Update/word_access_complete/$exit
      -- CP-element group 43: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_117_Update/word_access_complete/word_0/$exit
      -- CP-element group 43: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_117_Update/word_access_complete/word_0/ca
      -- CP-element group 43: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_117_Update/ptr_deref_117_Merge/$entry
      -- CP-element group 43: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_117_Update/ptr_deref_117_Merge/$exit
      -- CP-element group 43: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_117_Update/ptr_deref_117_Merge/merge_req
      -- CP-element group 43: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_117_Update/ptr_deref_117_Merge/merge_ack
      -- CP-element group 43: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_117_update_completed_
      -- 
    ca_603_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_117_load_0_ack_1, ack => maxPool4_CP_307_elements(43)); -- 
    -- CP-element group 44:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	28 
    -- CP-element group 44: marked-predecessors 
    -- CP-element group 44: 	46 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	46 
    -- CP-element group 44:  members (5) 
      -- CP-element group 44: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_121_sample_start_
      -- CP-element group 44: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_121_Sample/$entry
      -- CP-element group 44: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_121_Sample/word_access_start/$entry
      -- CP-element group 44: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_121_Sample/word_access_start/word_0/$entry
      -- CP-element group 44: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_121_Sample/word_access_start/word_0/rr
      -- 
    rr_641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(44), ack => ptr_deref_121_load_0_req_0); -- 
    maxPool4_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(28) & maxPool4_CP_307_elements(46);
      gj_maxPool4_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: marked-predecessors 
    -- CP-element group 45: 	47 
    -- CP-element group 45: 	182 
    -- CP-element group 45: 	186 
    -- CP-element group 45: 	190 
    -- CP-element group 45: 	194 
    -- CP-element group 45: 	198 
    -- CP-element group 45: 	202 
    -- CP-element group 45: 	206 
    -- CP-element group 45: 	210 
    -- CP-element group 45: 	214 
    -- CP-element group 45: 	218 
    -- CP-element group 45: 	222 
    -- CP-element group 45: 	226 
    -- CP-element group 45: 	230 
    -- CP-element group 45: 	234 
    -- CP-element group 45: 	238 
    -- CP-element group 45: 	242 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	47 
    -- CP-element group 45:  members (5) 
      -- CP-element group 45: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_121_update_start_
      -- CP-element group 45: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_121_Update/$entry
      -- CP-element group 45: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_121_Update/word_access_complete/$entry
      -- CP-element group 45: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_121_Update/word_access_complete/word_0/$entry
      -- CP-element group 45: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_121_Update/word_access_complete/word_0/cr
      -- 
    cr_652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(45), ack => ptr_deref_121_load_0_req_1); -- 
    maxPool4_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(47) & maxPool4_CP_307_elements(182) & maxPool4_CP_307_elements(186) & maxPool4_CP_307_elements(190) & maxPool4_CP_307_elements(194) & maxPool4_CP_307_elements(198) & maxPool4_CP_307_elements(202) & maxPool4_CP_307_elements(206) & maxPool4_CP_307_elements(210) & maxPool4_CP_307_elements(214) & maxPool4_CP_307_elements(218) & maxPool4_CP_307_elements(222) & maxPool4_CP_307_elements(226) & maxPool4_CP_307_elements(230) & maxPool4_CP_307_elements(234) & maxPool4_CP_307_elements(238) & maxPool4_CP_307_elements(242);
      gj_maxPool4_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	44 
    -- CP-element group 46: successors 
    -- CP-element group 46: marked-successors 
    -- CP-element group 46: 	23 
    -- CP-element group 46: 	44 
    -- CP-element group 46:  members (5) 
      -- CP-element group 46: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_121_sample_completed_
      -- CP-element group 46: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_121_Sample/$exit
      -- CP-element group 46: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_121_Sample/word_access_start/$exit
      -- CP-element group 46: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_121_Sample/word_access_start/word_0/$exit
      -- CP-element group 46: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_121_Sample/word_access_start/word_0/ra
      -- 
    ra_642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_121_load_0_ack_0, ack => maxPool4_CP_307_elements(46)); -- 
    -- CP-element group 47:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	45 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	180 
    -- CP-element group 47: 	184 
    -- CP-element group 47: 	188 
    -- CP-element group 47: 	192 
    -- CP-element group 47: 	196 
    -- CP-element group 47: 	200 
    -- CP-element group 47: 	204 
    -- CP-element group 47: 	208 
    -- CP-element group 47: 	212 
    -- CP-element group 47: 	216 
    -- CP-element group 47: 	220 
    -- CP-element group 47: 	224 
    -- CP-element group 47: 	228 
    -- CP-element group 47: 	232 
    -- CP-element group 47: 	236 
    -- CP-element group 47: 	240 
    -- CP-element group 47: marked-successors 
    -- CP-element group 47: 	45 
    -- CP-element group 47:  members (9) 
      -- CP-element group 47: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_121_update_completed_
      -- CP-element group 47: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_121_Update/$exit
      -- CP-element group 47: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_121_Update/word_access_complete/$exit
      -- CP-element group 47: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_121_Update/word_access_complete/word_0/$exit
      -- CP-element group 47: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_121_Update/word_access_complete/word_0/ca
      -- CP-element group 47: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_121_Update/ptr_deref_121_Merge/$entry
      -- CP-element group 47: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_121_Update/ptr_deref_121_Merge/$exit
      -- CP-element group 47: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_121_Update/ptr_deref_121_Merge/merge_req
      -- CP-element group 47: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_121_Update/ptr_deref_121_Merge/merge_ack
      -- 
    ca_653_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_121_load_0_ack_1, ack => maxPool4_CP_307_elements(47)); -- 
    -- CP-element group 48:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	35 
    -- CP-element group 48: marked-predecessors 
    -- CP-element group 48: 	50 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (5) 
      -- CP-element group 48: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_125_sample_start_
      -- CP-element group 48: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_125_Sample/$entry
      -- CP-element group 48: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_125_Sample/word_access_start/$entry
      -- CP-element group 48: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_125_Sample/word_access_start/word_0/$entry
      -- CP-element group 48: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_125_Sample/word_access_start/word_0/rr
      -- 
    rr_691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(48), ack => ptr_deref_125_load_0_req_0); -- 
    maxPool4_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(35) & maxPool4_CP_307_elements(50);
      gj_maxPool4_cp_element_group_48 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: marked-predecessors 
    -- CP-element group 49: 	51 
    -- CP-element group 49: 	246 
    -- CP-element group 49: 	250 
    -- CP-element group 49: 	254 
    -- CP-element group 49: 	258 
    -- CP-element group 49: 	262 
    -- CP-element group 49: 	266 
    -- CP-element group 49: 	270 
    -- CP-element group 49: 	274 
    -- CP-element group 49: 	278 
    -- CP-element group 49: 	282 
    -- CP-element group 49: 	286 
    -- CP-element group 49: 	290 
    -- CP-element group 49: 	294 
    -- CP-element group 49: 	298 
    -- CP-element group 49: 	302 
    -- CP-element group 49: 	306 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (5) 
      -- CP-element group 49: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_125_update_start_
      -- CP-element group 49: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_125_Update/$entry
      -- CP-element group 49: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_125_Update/word_access_complete/$entry
      -- CP-element group 49: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_125_Update/word_access_complete/word_0/$entry
      -- CP-element group 49: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_125_Update/word_access_complete/word_0/cr
      -- 
    cr_702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(49), ack => ptr_deref_125_load_0_req_1); -- 
    maxPool4_cp_element_group_49: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_49"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(51) & maxPool4_CP_307_elements(246) & maxPool4_CP_307_elements(250) & maxPool4_CP_307_elements(254) & maxPool4_CP_307_elements(258) & maxPool4_CP_307_elements(262) & maxPool4_CP_307_elements(266) & maxPool4_CP_307_elements(270) & maxPool4_CP_307_elements(274) & maxPool4_CP_307_elements(278) & maxPool4_CP_307_elements(282) & maxPool4_CP_307_elements(286) & maxPool4_CP_307_elements(290) & maxPool4_CP_307_elements(294) & maxPool4_CP_307_elements(298) & maxPool4_CP_307_elements(302) & maxPool4_CP_307_elements(306);
      gj_maxPool4_cp_element_group_49 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(49), clk => clk, reset => reset); --
    end block;
    -- CP-element group 50:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: successors 
    -- CP-element group 50: marked-successors 
    -- CP-element group 50: 	30 
    -- CP-element group 50: 	48 
    -- CP-element group 50:  members (5) 
      -- CP-element group 50: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_125_sample_completed_
      -- CP-element group 50: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_125_Sample/$exit
      -- CP-element group 50: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_125_Sample/word_access_start/$exit
      -- CP-element group 50: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_125_Sample/word_access_start/word_0/$exit
      -- CP-element group 50: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_125_Sample/word_access_start/word_0/ra
      -- 
    ra_692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_125_load_0_ack_0, ack => maxPool4_CP_307_elements(50)); -- 
    -- CP-element group 51:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	244 
    -- CP-element group 51: 	248 
    -- CP-element group 51: 	252 
    -- CP-element group 51: 	256 
    -- CP-element group 51: 	260 
    -- CP-element group 51: 	264 
    -- CP-element group 51: 	268 
    -- CP-element group 51: 	272 
    -- CP-element group 51: 	276 
    -- CP-element group 51: 	280 
    -- CP-element group 51: 	284 
    -- CP-element group 51: 	288 
    -- CP-element group 51: 	292 
    -- CP-element group 51: 	296 
    -- CP-element group 51: 	300 
    -- CP-element group 51: 	304 
    -- CP-element group 51: marked-successors 
    -- CP-element group 51: 	49 
    -- CP-element group 51:  members (9) 
      -- CP-element group 51: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_125_update_completed_
      -- CP-element group 51: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_125_Update/$exit
      -- CP-element group 51: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_125_Update/word_access_complete/$exit
      -- CP-element group 51: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_125_Update/word_access_complete/word_0/$exit
      -- CP-element group 51: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_125_Update/word_access_complete/word_0/ca
      -- CP-element group 51: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_125_Update/ptr_deref_125_Merge/$entry
      -- CP-element group 51: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_125_Update/ptr_deref_125_Merge/$exit
      -- CP-element group 51: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_125_Update/ptr_deref_125_Merge/merge_req
      -- CP-element group 51: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_125_Update/ptr_deref_125_Merge/merge_ack
      -- 
    ca_703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_125_load_0_ack_1, ack => maxPool4_CP_307_elements(51)); -- 
    -- CP-element group 52:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	39 
    -- CP-element group 52: marked-predecessors 
    -- CP-element group 52: 	54 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 assign_stmt_89_to_assign_stmt_1130/slice_130_sample_start_
      -- CP-element group 52: 	 assign_stmt_89_to_assign_stmt_1130/slice_130_Sample/$entry
      -- CP-element group 52: 	 assign_stmt_89_to_assign_stmt_1130/slice_130_Sample/rr
      -- 
    rr_716_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_716_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(52), ack => slice_130_inst_req_0); -- 
    maxPool4_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(39) & maxPool4_CP_307_elements(54);
      gj_maxPool4_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: marked-predecessors 
    -- CP-element group 53: 	55 
    -- CP-element group 53: 	321 
    -- CP-element group 53: 	386 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 assign_stmt_89_to_assign_stmt_1130/slice_130_update_start_
      -- CP-element group 53: 	 assign_stmt_89_to_assign_stmt_1130/slice_130_Update/$entry
      -- CP-element group 53: 	 assign_stmt_89_to_assign_stmt_1130/slice_130_Update/cr
      -- 
    cr_721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(53), ack => slice_130_inst_req_1); -- 
    maxPool4_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(55) & maxPool4_CP_307_elements(321) & maxPool4_CP_307_elements(386);
      gj_maxPool4_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: marked-successors 
    -- CP-element group 54: 	37 
    -- CP-element group 54: 	52 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 assign_stmt_89_to_assign_stmt_1130/slice_130_sample_completed_
      -- CP-element group 54: 	 assign_stmt_89_to_assign_stmt_1130/slice_130_Sample/$exit
      -- CP-element group 54: 	 assign_stmt_89_to_assign_stmt_1130/slice_130_Sample/ra
      -- 
    ra_717_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_130_inst_ack_0, ack => maxPool4_CP_307_elements(54)); -- 
    -- CP-element group 55:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	319 
    -- CP-element group 55: 	384 
    -- CP-element group 55: marked-successors 
    -- CP-element group 55: 	53 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 assign_stmt_89_to_assign_stmt_1130/slice_130_update_completed_
      -- CP-element group 55: 	 assign_stmt_89_to_assign_stmt_1130/slice_130_Update/$exit
      -- CP-element group 55: 	 assign_stmt_89_to_assign_stmt_1130/slice_130_Update/ca
      -- 
    ca_722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_130_inst_ack_1, ack => maxPool4_CP_307_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	39 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	58 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 assign_stmt_89_to_assign_stmt_1130/slice_134_sample_start_
      -- CP-element group 56: 	 assign_stmt_89_to_assign_stmt_1130/slice_134_Sample/$entry
      -- CP-element group 56: 	 assign_stmt_89_to_assign_stmt_1130/slice_134_Sample/rr
      -- 
    rr_730_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_730_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(56), ack => slice_134_inst_req_0); -- 
    maxPool4_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(39) & maxPool4_CP_307_elements(58);
      gj_maxPool4_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: marked-predecessors 
    -- CP-element group 57: 	59 
    -- CP-element group 57: 	321 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 assign_stmt_89_to_assign_stmt_1130/slice_134_update_start_
      -- CP-element group 57: 	 assign_stmt_89_to_assign_stmt_1130/slice_134_Update/$entry
      -- CP-element group 57: 	 assign_stmt_89_to_assign_stmt_1130/slice_134_Update/cr
      -- 
    cr_735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(57), ack => slice_134_inst_req_1); -- 
    maxPool4_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(59) & maxPool4_CP_307_elements(321);
      gj_maxPool4_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58: marked-successors 
    -- CP-element group 58: 	37 
    -- CP-element group 58: 	56 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 assign_stmt_89_to_assign_stmt_1130/slice_134_sample_completed_
      -- CP-element group 58: 	 assign_stmt_89_to_assign_stmt_1130/slice_134_Sample/$exit
      -- CP-element group 58: 	 assign_stmt_89_to_assign_stmt_1130/slice_134_Sample/ra
      -- 
    ra_731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_134_inst_ack_0, ack => maxPool4_CP_307_elements(58)); -- 
    -- CP-element group 59:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	319 
    -- CP-element group 59: marked-successors 
    -- CP-element group 59: 	57 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 assign_stmt_89_to_assign_stmt_1130/slice_134_update_completed_
      -- CP-element group 59: 	 assign_stmt_89_to_assign_stmt_1130/slice_134_Update/$exit
      -- CP-element group 59: 	 assign_stmt_89_to_assign_stmt_1130/slice_134_Update/ca
      -- 
    ca_736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_134_inst_ack_1, ack => maxPool4_CP_307_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	39 
    -- CP-element group 60: marked-predecessors 
    -- CP-element group 60: 	62 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 assign_stmt_89_to_assign_stmt_1130/slice_138_sample_start_
      -- CP-element group 60: 	 assign_stmt_89_to_assign_stmt_1130/slice_138_Sample/$entry
      -- CP-element group 60: 	 assign_stmt_89_to_assign_stmt_1130/slice_138_Sample/rr
      -- 
    rr_744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(60), ack => slice_138_inst_req_0); -- 
    maxPool4_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(39) & maxPool4_CP_307_elements(62);
      gj_maxPool4_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: marked-predecessors 
    -- CP-element group 61: 	63 
    -- CP-element group 61: 	321 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 assign_stmt_89_to_assign_stmt_1130/slice_138_update_start_
      -- CP-element group 61: 	 assign_stmt_89_to_assign_stmt_1130/slice_138_Update/$entry
      -- CP-element group 61: 	 assign_stmt_89_to_assign_stmt_1130/slice_138_Update/cr
      -- 
    cr_749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(61), ack => slice_138_inst_req_1); -- 
    maxPool4_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(63) & maxPool4_CP_307_elements(321);
      gj_maxPool4_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: marked-successors 
    -- CP-element group 62: 	37 
    -- CP-element group 62: 	60 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 assign_stmt_89_to_assign_stmt_1130/slice_138_sample_completed_
      -- CP-element group 62: 	 assign_stmt_89_to_assign_stmt_1130/slice_138_Sample/$exit
      -- CP-element group 62: 	 assign_stmt_89_to_assign_stmt_1130/slice_138_Sample/ra
      -- 
    ra_745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_138_inst_ack_0, ack => maxPool4_CP_307_elements(62)); -- 
    -- CP-element group 63:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	319 
    -- CP-element group 63: marked-successors 
    -- CP-element group 63: 	61 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 assign_stmt_89_to_assign_stmt_1130/slice_138_update_completed_
      -- CP-element group 63: 	 assign_stmt_89_to_assign_stmt_1130/slice_138_Update/$exit
      -- CP-element group 63: 	 assign_stmt_89_to_assign_stmt_1130/slice_138_Update/ca
      -- 
    ca_750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_138_inst_ack_1, ack => maxPool4_CP_307_elements(63)); -- 
    -- CP-element group 64:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	39 
    -- CP-element group 64: marked-predecessors 
    -- CP-element group 64: 	66 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 assign_stmt_89_to_assign_stmt_1130/slice_142_sample_start_
      -- CP-element group 64: 	 assign_stmt_89_to_assign_stmt_1130/slice_142_Sample/$entry
      -- CP-element group 64: 	 assign_stmt_89_to_assign_stmt_1130/slice_142_Sample/rr
      -- 
    rr_758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(64), ack => slice_142_inst_req_0); -- 
    maxPool4_cp_element_group_64: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_64"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(39) & maxPool4_CP_307_elements(66);
      gj_maxPool4_cp_element_group_64 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(64), clk => clk, reset => reset); --
    end block;
    -- CP-element group 65:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: marked-predecessors 
    -- CP-element group 65: 	67 
    -- CP-element group 65: 	321 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 assign_stmt_89_to_assign_stmt_1130/slice_142_update_start_
      -- CP-element group 65: 	 assign_stmt_89_to_assign_stmt_1130/slice_142_Update/$entry
      -- CP-element group 65: 	 assign_stmt_89_to_assign_stmt_1130/slice_142_Update/cr
      -- 
    cr_763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(65), ack => slice_142_inst_req_1); -- 
    maxPool4_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(67) & maxPool4_CP_307_elements(321);
      gj_maxPool4_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66: marked-successors 
    -- CP-element group 66: 	37 
    -- CP-element group 66: 	64 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 assign_stmt_89_to_assign_stmt_1130/slice_142_sample_completed_
      -- CP-element group 66: 	 assign_stmt_89_to_assign_stmt_1130/slice_142_Sample/$exit
      -- CP-element group 66: 	 assign_stmt_89_to_assign_stmt_1130/slice_142_Sample/ra
      -- 
    ra_759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_142_inst_ack_0, ack => maxPool4_CP_307_elements(66)); -- 
    -- CP-element group 67:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	319 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	65 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 assign_stmt_89_to_assign_stmt_1130/slice_142_update_completed_
      -- CP-element group 67: 	 assign_stmt_89_to_assign_stmt_1130/slice_142_Update/$exit
      -- CP-element group 67: 	 assign_stmt_89_to_assign_stmt_1130/slice_142_Update/ca
      -- 
    ca_764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_142_inst_ack_1, ack => maxPool4_CP_307_elements(67)); -- 
    -- CP-element group 68:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	39 
    -- CP-element group 68: marked-predecessors 
    -- CP-element group 68: 	70 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 assign_stmt_89_to_assign_stmt_1130/slice_146_sample_start_
      -- CP-element group 68: 	 assign_stmt_89_to_assign_stmt_1130/slice_146_Sample/$entry
      -- CP-element group 68: 	 assign_stmt_89_to_assign_stmt_1130/slice_146_Sample/rr
      -- 
    rr_772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(68), ack => slice_146_inst_req_0); -- 
    maxPool4_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(39) & maxPool4_CP_307_elements(70);
      gj_maxPool4_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: marked-predecessors 
    -- CP-element group 69: 	71 
    -- CP-element group 69: 	340 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 assign_stmt_89_to_assign_stmt_1130/slice_146_update_start_
      -- CP-element group 69: 	 assign_stmt_89_to_assign_stmt_1130/slice_146_Update/$entry
      -- CP-element group 69: 	 assign_stmt_89_to_assign_stmt_1130/slice_146_Update/cr
      -- 
    cr_777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(69), ack => slice_146_inst_req_1); -- 
    maxPool4_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(71) & maxPool4_CP_307_elements(340);
      gj_maxPool4_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: marked-successors 
    -- CP-element group 70: 	37 
    -- CP-element group 70: 	68 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 assign_stmt_89_to_assign_stmt_1130/slice_146_sample_completed_
      -- CP-element group 70: 	 assign_stmt_89_to_assign_stmt_1130/slice_146_Sample/$exit
      -- CP-element group 70: 	 assign_stmt_89_to_assign_stmt_1130/slice_146_Sample/ra
      -- 
    ra_773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_146_inst_ack_0, ack => maxPool4_CP_307_elements(70)); -- 
    -- CP-element group 71:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	338 
    -- CP-element group 71: marked-successors 
    -- CP-element group 71: 	69 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 assign_stmt_89_to_assign_stmt_1130/slice_146_update_completed_
      -- CP-element group 71: 	 assign_stmt_89_to_assign_stmt_1130/slice_146_Update/$exit
      -- CP-element group 71: 	 assign_stmt_89_to_assign_stmt_1130/slice_146_Update/ca
      -- 
    ca_778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_146_inst_ack_1, ack => maxPool4_CP_307_elements(71)); -- 
    -- CP-element group 72:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	39 
    -- CP-element group 72: marked-predecessors 
    -- CP-element group 72: 	74 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 assign_stmt_89_to_assign_stmt_1130/slice_150_sample_start_
      -- CP-element group 72: 	 assign_stmt_89_to_assign_stmt_1130/slice_150_Sample/$entry
      -- CP-element group 72: 	 assign_stmt_89_to_assign_stmt_1130/slice_150_Sample/rr
      -- 
    rr_786_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_786_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(72), ack => slice_150_inst_req_0); -- 
    maxPool4_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(39) & maxPool4_CP_307_elements(74);
      gj_maxPool4_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: marked-predecessors 
    -- CP-element group 73: 	75 
    -- CP-element group 73: 	340 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 assign_stmt_89_to_assign_stmt_1130/slice_150_update_start_
      -- CP-element group 73: 	 assign_stmt_89_to_assign_stmt_1130/slice_150_Update/$entry
      -- CP-element group 73: 	 assign_stmt_89_to_assign_stmt_1130/slice_150_Update/cr
      -- 
    cr_791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(73), ack => slice_150_inst_req_1); -- 
    maxPool4_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(75) & maxPool4_CP_307_elements(340);
      gj_maxPool4_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: successors 
    -- CP-element group 74: marked-successors 
    -- CP-element group 74: 	37 
    -- CP-element group 74: 	72 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 assign_stmt_89_to_assign_stmt_1130/slice_150_sample_completed_
      -- CP-element group 74: 	 assign_stmt_89_to_assign_stmt_1130/slice_150_Sample/$exit
      -- CP-element group 74: 	 assign_stmt_89_to_assign_stmt_1130/slice_150_Sample/ra
      -- 
    ra_787_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_150_inst_ack_0, ack => maxPool4_CP_307_elements(74)); -- 
    -- CP-element group 75:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	338 
    -- CP-element group 75: marked-successors 
    -- CP-element group 75: 	73 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 assign_stmt_89_to_assign_stmt_1130/slice_150_update_completed_
      -- CP-element group 75: 	 assign_stmt_89_to_assign_stmt_1130/slice_150_Update/$exit
      -- CP-element group 75: 	 assign_stmt_89_to_assign_stmt_1130/slice_150_Update/ca
      -- 
    ca_792_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_150_inst_ack_1, ack => maxPool4_CP_307_elements(75)); -- 
    -- CP-element group 76:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	39 
    -- CP-element group 76: marked-predecessors 
    -- CP-element group 76: 	78 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 assign_stmt_89_to_assign_stmt_1130/slice_154_sample_start_
      -- CP-element group 76: 	 assign_stmt_89_to_assign_stmt_1130/slice_154_Sample/$entry
      -- CP-element group 76: 	 assign_stmt_89_to_assign_stmt_1130/slice_154_Sample/rr
      -- 
    rr_800_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_800_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(76), ack => slice_154_inst_req_0); -- 
    maxPool4_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(39) & maxPool4_CP_307_elements(78);
      gj_maxPool4_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: marked-predecessors 
    -- CP-element group 77: 	79 
    -- CP-element group 77: 	340 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	79 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 assign_stmt_89_to_assign_stmt_1130/slice_154_update_start_
      -- CP-element group 77: 	 assign_stmt_89_to_assign_stmt_1130/slice_154_Update/$entry
      -- CP-element group 77: 	 assign_stmt_89_to_assign_stmt_1130/slice_154_Update/cr
      -- 
    cr_805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(77), ack => slice_154_inst_req_1); -- 
    maxPool4_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(79) & maxPool4_CP_307_elements(340);
      gj_maxPool4_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: successors 
    -- CP-element group 78: marked-successors 
    -- CP-element group 78: 	37 
    -- CP-element group 78: 	76 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 assign_stmt_89_to_assign_stmt_1130/slice_154_sample_completed_
      -- CP-element group 78: 	 assign_stmt_89_to_assign_stmt_1130/slice_154_Sample/$exit
      -- CP-element group 78: 	 assign_stmt_89_to_assign_stmt_1130/slice_154_Sample/ra
      -- 
    ra_801_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_154_inst_ack_0, ack => maxPool4_CP_307_elements(78)); -- 
    -- CP-element group 79:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	338 
    -- CP-element group 79: marked-successors 
    -- CP-element group 79: 	77 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 assign_stmt_89_to_assign_stmt_1130/slice_154_update_completed_
      -- CP-element group 79: 	 assign_stmt_89_to_assign_stmt_1130/slice_154_Update/$exit
      -- CP-element group 79: 	 assign_stmt_89_to_assign_stmt_1130/slice_154_Update/ca
      -- 
    ca_806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_154_inst_ack_1, ack => maxPool4_CP_307_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	39 
    -- CP-element group 80: marked-predecessors 
    -- CP-element group 80: 	82 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 assign_stmt_89_to_assign_stmt_1130/slice_158_sample_start_
      -- CP-element group 80: 	 assign_stmt_89_to_assign_stmt_1130/slice_158_Sample/$entry
      -- CP-element group 80: 	 assign_stmt_89_to_assign_stmt_1130/slice_158_Sample/rr
      -- 
    rr_814_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_814_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(80), ack => slice_158_inst_req_0); -- 
    maxPool4_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(39) & maxPool4_CP_307_elements(82);
      gj_maxPool4_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: marked-predecessors 
    -- CP-element group 81: 	83 
    -- CP-element group 81: 	340 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 assign_stmt_89_to_assign_stmt_1130/slice_158_update_start_
      -- CP-element group 81: 	 assign_stmt_89_to_assign_stmt_1130/slice_158_Update/$entry
      -- CP-element group 81: 	 assign_stmt_89_to_assign_stmt_1130/slice_158_Update/cr
      -- 
    cr_819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(81), ack => slice_158_inst_req_1); -- 
    maxPool4_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(83) & maxPool4_CP_307_elements(340);
      gj_maxPool4_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: successors 
    -- CP-element group 82: marked-successors 
    -- CP-element group 82: 	37 
    -- CP-element group 82: 	80 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 assign_stmt_89_to_assign_stmt_1130/slice_158_sample_completed_
      -- CP-element group 82: 	 assign_stmt_89_to_assign_stmt_1130/slice_158_Sample/$exit
      -- CP-element group 82: 	 assign_stmt_89_to_assign_stmt_1130/slice_158_Sample/ra
      -- 
    ra_815_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_158_inst_ack_0, ack => maxPool4_CP_307_elements(82)); -- 
    -- CP-element group 83:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	338 
    -- CP-element group 83: marked-successors 
    -- CP-element group 83: 	81 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 assign_stmt_89_to_assign_stmt_1130/slice_158_update_completed_
      -- CP-element group 83: 	 assign_stmt_89_to_assign_stmt_1130/slice_158_Update/$exit
      -- CP-element group 83: 	 assign_stmt_89_to_assign_stmt_1130/slice_158_Update/ca
      -- 
    ca_820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_158_inst_ack_1, ack => maxPool4_CP_307_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	39 
    -- CP-element group 84: marked-predecessors 
    -- CP-element group 84: 	86 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 assign_stmt_89_to_assign_stmt_1130/slice_162_sample_start_
      -- CP-element group 84: 	 assign_stmt_89_to_assign_stmt_1130/slice_162_Sample/$entry
      -- CP-element group 84: 	 assign_stmt_89_to_assign_stmt_1130/slice_162_Sample/rr
      -- 
    rr_828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(84), ack => slice_162_inst_req_0); -- 
    maxPool4_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(39) & maxPool4_CP_307_elements(86);
      gj_maxPool4_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: marked-predecessors 
    -- CP-element group 85: 	87 
    -- CP-element group 85: 	359 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 assign_stmt_89_to_assign_stmt_1130/slice_162_update_start_
      -- CP-element group 85: 	 assign_stmt_89_to_assign_stmt_1130/slice_162_Update/$entry
      -- CP-element group 85: 	 assign_stmt_89_to_assign_stmt_1130/slice_162_Update/cr
      -- 
    cr_833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(85), ack => slice_162_inst_req_1); -- 
    maxPool4_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(87) & maxPool4_CP_307_elements(359);
      gj_maxPool4_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: successors 
    -- CP-element group 86: marked-successors 
    -- CP-element group 86: 	37 
    -- CP-element group 86: 	84 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 assign_stmt_89_to_assign_stmt_1130/slice_162_sample_completed_
      -- CP-element group 86: 	 assign_stmt_89_to_assign_stmt_1130/slice_162_Sample/$exit
      -- CP-element group 86: 	 assign_stmt_89_to_assign_stmt_1130/slice_162_Sample/ra
      -- 
    ra_829_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_162_inst_ack_0, ack => maxPool4_CP_307_elements(86)); -- 
    -- CP-element group 87:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	357 
    -- CP-element group 87: marked-successors 
    -- CP-element group 87: 	85 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 assign_stmt_89_to_assign_stmt_1130/slice_162_update_completed_
      -- CP-element group 87: 	 assign_stmt_89_to_assign_stmt_1130/slice_162_Update/$exit
      -- CP-element group 87: 	 assign_stmt_89_to_assign_stmt_1130/slice_162_Update/ca
      -- 
    ca_834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_162_inst_ack_1, ack => maxPool4_CP_307_elements(87)); -- 
    -- CP-element group 88:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	39 
    -- CP-element group 88: marked-predecessors 
    -- CP-element group 88: 	90 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 assign_stmt_89_to_assign_stmt_1130/slice_166_sample_start_
      -- CP-element group 88: 	 assign_stmt_89_to_assign_stmt_1130/slice_166_Sample/$entry
      -- CP-element group 88: 	 assign_stmt_89_to_assign_stmt_1130/slice_166_Sample/rr
      -- 
    rr_842_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_842_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(88), ack => slice_166_inst_req_0); -- 
    maxPool4_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(39) & maxPool4_CP_307_elements(90);
      gj_maxPool4_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: marked-predecessors 
    -- CP-element group 89: 	91 
    -- CP-element group 89: 	359 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 assign_stmt_89_to_assign_stmt_1130/slice_166_update_start_
      -- CP-element group 89: 	 assign_stmt_89_to_assign_stmt_1130/slice_166_Update/$entry
      -- CP-element group 89: 	 assign_stmt_89_to_assign_stmt_1130/slice_166_Update/cr
      -- 
    cr_847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(89), ack => slice_166_inst_req_1); -- 
    maxPool4_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(91) & maxPool4_CP_307_elements(359);
      gj_maxPool4_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: successors 
    -- CP-element group 90: marked-successors 
    -- CP-element group 90: 	37 
    -- CP-element group 90: 	88 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 assign_stmt_89_to_assign_stmt_1130/slice_166_sample_completed_
      -- CP-element group 90: 	 assign_stmt_89_to_assign_stmt_1130/slice_166_Sample/$exit
      -- CP-element group 90: 	 assign_stmt_89_to_assign_stmt_1130/slice_166_Sample/ra
      -- 
    ra_843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_166_inst_ack_0, ack => maxPool4_CP_307_elements(90)); -- 
    -- CP-element group 91:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	357 
    -- CP-element group 91: marked-successors 
    -- CP-element group 91: 	89 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 assign_stmt_89_to_assign_stmt_1130/slice_166_update_completed_
      -- CP-element group 91: 	 assign_stmt_89_to_assign_stmt_1130/slice_166_Update/$exit
      -- CP-element group 91: 	 assign_stmt_89_to_assign_stmt_1130/slice_166_Update/ca
      -- 
    ca_848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_166_inst_ack_1, ack => maxPool4_CP_307_elements(91)); -- 
    -- CP-element group 92:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	39 
    -- CP-element group 92: marked-predecessors 
    -- CP-element group 92: 	94 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 assign_stmt_89_to_assign_stmt_1130/slice_170_sample_start_
      -- CP-element group 92: 	 assign_stmt_89_to_assign_stmt_1130/slice_170_Sample/$entry
      -- CP-element group 92: 	 assign_stmt_89_to_assign_stmt_1130/slice_170_Sample/rr
      -- 
    rr_856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(92), ack => slice_170_inst_req_0); -- 
    maxPool4_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(39) & maxPool4_CP_307_elements(94);
      gj_maxPool4_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: marked-predecessors 
    -- CP-element group 93: 	95 
    -- CP-element group 93: 	359 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 assign_stmt_89_to_assign_stmt_1130/slice_170_update_start_
      -- CP-element group 93: 	 assign_stmt_89_to_assign_stmt_1130/slice_170_Update/$entry
      -- CP-element group 93: 	 assign_stmt_89_to_assign_stmt_1130/slice_170_Update/cr
      -- 
    cr_861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(93), ack => slice_170_inst_req_1); -- 
    maxPool4_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(95) & maxPool4_CP_307_elements(359);
      gj_maxPool4_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: successors 
    -- CP-element group 94: marked-successors 
    -- CP-element group 94: 	37 
    -- CP-element group 94: 	92 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 assign_stmt_89_to_assign_stmt_1130/slice_170_sample_completed_
      -- CP-element group 94: 	 assign_stmt_89_to_assign_stmt_1130/slice_170_Sample/$exit
      -- CP-element group 94: 	 assign_stmt_89_to_assign_stmt_1130/slice_170_Sample/ra
      -- 
    ra_857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_170_inst_ack_0, ack => maxPool4_CP_307_elements(94)); -- 
    -- CP-element group 95:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	357 
    -- CP-element group 95: marked-successors 
    -- CP-element group 95: 	93 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 assign_stmt_89_to_assign_stmt_1130/slice_170_update_completed_
      -- CP-element group 95: 	 assign_stmt_89_to_assign_stmt_1130/slice_170_Update/$exit
      -- CP-element group 95: 	 assign_stmt_89_to_assign_stmt_1130/slice_170_Update/ca
      -- 
    ca_862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_170_inst_ack_1, ack => maxPool4_CP_307_elements(95)); -- 
    -- CP-element group 96:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	39 
    -- CP-element group 96: marked-predecessors 
    -- CP-element group 96: 	98 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	98 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 assign_stmt_89_to_assign_stmt_1130/slice_174_sample_start_
      -- CP-element group 96: 	 assign_stmt_89_to_assign_stmt_1130/slice_174_Sample/$entry
      -- CP-element group 96: 	 assign_stmt_89_to_assign_stmt_1130/slice_174_Sample/rr
      -- 
    rr_870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(96), ack => slice_174_inst_req_0); -- 
    maxPool4_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(39) & maxPool4_CP_307_elements(98);
      gj_maxPool4_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: marked-predecessors 
    -- CP-element group 97: 	99 
    -- CP-element group 97: 	359 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	99 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 assign_stmt_89_to_assign_stmt_1130/slice_174_update_start_
      -- CP-element group 97: 	 assign_stmt_89_to_assign_stmt_1130/slice_174_Update/$entry
      -- CP-element group 97: 	 assign_stmt_89_to_assign_stmt_1130/slice_174_Update/cr
      -- 
    cr_875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(97), ack => slice_174_inst_req_1); -- 
    maxPool4_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(99) & maxPool4_CP_307_elements(359);
      gj_maxPool4_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	96 
    -- CP-element group 98: successors 
    -- CP-element group 98: marked-successors 
    -- CP-element group 98: 	37 
    -- CP-element group 98: 	96 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 assign_stmt_89_to_assign_stmt_1130/slice_174_sample_completed_
      -- CP-element group 98: 	 assign_stmt_89_to_assign_stmt_1130/slice_174_Sample/$exit
      -- CP-element group 98: 	 assign_stmt_89_to_assign_stmt_1130/slice_174_Sample/ra
      -- 
    ra_871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_174_inst_ack_0, ack => maxPool4_CP_307_elements(98)); -- 
    -- CP-element group 99:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	97 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	357 
    -- CP-element group 99: marked-successors 
    -- CP-element group 99: 	97 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 assign_stmt_89_to_assign_stmt_1130/slice_174_update_completed_
      -- CP-element group 99: 	 assign_stmt_89_to_assign_stmt_1130/slice_174_Update/$exit
      -- CP-element group 99: 	 assign_stmt_89_to_assign_stmt_1130/slice_174_Update/ca
      -- 
    ca_876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_174_inst_ack_1, ack => maxPool4_CP_307_elements(99)); -- 
    -- CP-element group 100:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	39 
    -- CP-element group 100: marked-predecessors 
    -- CP-element group 100: 	102 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	102 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 assign_stmt_89_to_assign_stmt_1130/slice_178_sample_start_
      -- CP-element group 100: 	 assign_stmt_89_to_assign_stmt_1130/slice_178_Sample/$entry
      -- CP-element group 100: 	 assign_stmt_89_to_assign_stmt_1130/slice_178_Sample/rr
      -- 
    rr_884_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_884_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(100), ack => slice_178_inst_req_0); -- 
    maxPool4_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(39) & maxPool4_CP_307_elements(102);
      gj_maxPool4_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: marked-predecessors 
    -- CP-element group 101: 	103 
    -- CP-element group 101: 	378 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	103 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 assign_stmt_89_to_assign_stmt_1130/slice_178_update_start_
      -- CP-element group 101: 	 assign_stmt_89_to_assign_stmt_1130/slice_178_Update/$entry
      -- CP-element group 101: 	 assign_stmt_89_to_assign_stmt_1130/slice_178_Update/cr
      -- 
    cr_889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(101), ack => slice_178_inst_req_1); -- 
    maxPool4_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(103) & maxPool4_CP_307_elements(378);
      gj_maxPool4_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	100 
    -- CP-element group 102: successors 
    -- CP-element group 102: marked-successors 
    -- CP-element group 102: 	37 
    -- CP-element group 102: 	100 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 assign_stmt_89_to_assign_stmt_1130/slice_178_sample_completed_
      -- CP-element group 102: 	 assign_stmt_89_to_assign_stmt_1130/slice_178_Sample/$exit
      -- CP-element group 102: 	 assign_stmt_89_to_assign_stmt_1130/slice_178_Sample/ra
      -- 
    ra_885_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_178_inst_ack_0, ack => maxPool4_CP_307_elements(102)); -- 
    -- CP-element group 103:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	376 
    -- CP-element group 103: marked-successors 
    -- CP-element group 103: 	101 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 assign_stmt_89_to_assign_stmt_1130/slice_178_update_completed_
      -- CP-element group 103: 	 assign_stmt_89_to_assign_stmt_1130/slice_178_Update/$exit
      -- CP-element group 103: 	 assign_stmt_89_to_assign_stmt_1130/slice_178_Update/ca
      -- 
    ca_890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_178_inst_ack_1, ack => maxPool4_CP_307_elements(103)); -- 
    -- CP-element group 104:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	39 
    -- CP-element group 104: marked-predecessors 
    -- CP-element group 104: 	106 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	106 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 assign_stmt_89_to_assign_stmt_1130/slice_182_sample_start_
      -- CP-element group 104: 	 assign_stmt_89_to_assign_stmt_1130/slice_182_Sample/$entry
      -- CP-element group 104: 	 assign_stmt_89_to_assign_stmt_1130/slice_182_Sample/rr
      -- 
    rr_898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(104), ack => slice_182_inst_req_0); -- 
    maxPool4_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(39) & maxPool4_CP_307_elements(106);
      gj_maxPool4_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: marked-predecessors 
    -- CP-element group 105: 	107 
    -- CP-element group 105: 	378 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 assign_stmt_89_to_assign_stmt_1130/slice_182_update_start_
      -- CP-element group 105: 	 assign_stmt_89_to_assign_stmt_1130/slice_182_Update/$entry
      -- CP-element group 105: 	 assign_stmt_89_to_assign_stmt_1130/slice_182_Update/cr
      -- 
    cr_903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(105), ack => slice_182_inst_req_1); -- 
    maxPool4_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(107) & maxPool4_CP_307_elements(378);
      gj_maxPool4_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	104 
    -- CP-element group 106: successors 
    -- CP-element group 106: marked-successors 
    -- CP-element group 106: 	37 
    -- CP-element group 106: 	104 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 assign_stmt_89_to_assign_stmt_1130/slice_182_sample_completed_
      -- CP-element group 106: 	 assign_stmt_89_to_assign_stmt_1130/slice_182_Sample/$exit
      -- CP-element group 106: 	 assign_stmt_89_to_assign_stmt_1130/slice_182_Sample/ra
      -- 
    ra_899_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_182_inst_ack_0, ack => maxPool4_CP_307_elements(106)); -- 
    -- CP-element group 107:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	376 
    -- CP-element group 107: marked-successors 
    -- CP-element group 107: 	105 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 assign_stmt_89_to_assign_stmt_1130/slice_182_update_completed_
      -- CP-element group 107: 	 assign_stmt_89_to_assign_stmt_1130/slice_182_Update/$exit
      -- CP-element group 107: 	 assign_stmt_89_to_assign_stmt_1130/slice_182_Update/ca
      -- 
    ca_904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_182_inst_ack_1, ack => maxPool4_CP_307_elements(107)); -- 
    -- CP-element group 108:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	39 
    -- CP-element group 108: marked-predecessors 
    -- CP-element group 108: 	110 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	110 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 assign_stmt_89_to_assign_stmt_1130/slice_186_sample_start_
      -- CP-element group 108: 	 assign_stmt_89_to_assign_stmt_1130/slice_186_Sample/$entry
      -- CP-element group 108: 	 assign_stmt_89_to_assign_stmt_1130/slice_186_Sample/rr
      -- 
    rr_912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(108), ack => slice_186_inst_req_0); -- 
    maxPool4_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(39) & maxPool4_CP_307_elements(110);
      gj_maxPool4_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: marked-predecessors 
    -- CP-element group 109: 	111 
    -- CP-element group 109: 	378 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 assign_stmt_89_to_assign_stmt_1130/slice_186_update_start_
      -- CP-element group 109: 	 assign_stmt_89_to_assign_stmt_1130/slice_186_Update/$entry
      -- CP-element group 109: 	 assign_stmt_89_to_assign_stmt_1130/slice_186_Update/cr
      -- 
    cr_917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(109), ack => slice_186_inst_req_1); -- 
    maxPool4_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(111) & maxPool4_CP_307_elements(378);
      gj_maxPool4_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	108 
    -- CP-element group 110: successors 
    -- CP-element group 110: marked-successors 
    -- CP-element group 110: 	37 
    -- CP-element group 110: 	108 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 assign_stmt_89_to_assign_stmt_1130/slice_186_sample_completed_
      -- CP-element group 110: 	 assign_stmt_89_to_assign_stmt_1130/slice_186_Sample/$exit
      -- CP-element group 110: 	 assign_stmt_89_to_assign_stmt_1130/slice_186_Sample/ra
      -- 
    ra_913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_186_inst_ack_0, ack => maxPool4_CP_307_elements(110)); -- 
    -- CP-element group 111:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	376 
    -- CP-element group 111: marked-successors 
    -- CP-element group 111: 	109 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 assign_stmt_89_to_assign_stmt_1130/slice_186_update_completed_
      -- CP-element group 111: 	 assign_stmt_89_to_assign_stmt_1130/slice_186_Update/$exit
      -- CP-element group 111: 	 assign_stmt_89_to_assign_stmt_1130/slice_186_Update/ca
      -- 
    ca_918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_186_inst_ack_1, ack => maxPool4_CP_307_elements(111)); -- 
    -- CP-element group 112:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	39 
    -- CP-element group 112: marked-predecessors 
    -- CP-element group 112: 	114 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 assign_stmt_89_to_assign_stmt_1130/slice_190_sample_start_
      -- CP-element group 112: 	 assign_stmt_89_to_assign_stmt_1130/slice_190_Sample/$entry
      -- CP-element group 112: 	 assign_stmt_89_to_assign_stmt_1130/slice_190_Sample/rr
      -- 
    rr_926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(112), ack => slice_190_inst_req_0); -- 
    maxPool4_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(39) & maxPool4_CP_307_elements(114);
      gj_maxPool4_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: marked-predecessors 
    -- CP-element group 113: 	115 
    -- CP-element group 113: 	378 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 assign_stmt_89_to_assign_stmt_1130/slice_190_update_start_
      -- CP-element group 113: 	 assign_stmt_89_to_assign_stmt_1130/slice_190_Update/$entry
      -- CP-element group 113: 	 assign_stmt_89_to_assign_stmt_1130/slice_190_Update/cr
      -- 
    cr_931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(113), ack => slice_190_inst_req_1); -- 
    maxPool4_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(115) & maxPool4_CP_307_elements(378);
      gj_maxPool4_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: successors 
    -- CP-element group 114: marked-successors 
    -- CP-element group 114: 	37 
    -- CP-element group 114: 	112 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 assign_stmt_89_to_assign_stmt_1130/slice_190_sample_completed_
      -- CP-element group 114: 	 assign_stmt_89_to_assign_stmt_1130/slice_190_Sample/$exit
      -- CP-element group 114: 	 assign_stmt_89_to_assign_stmt_1130/slice_190_Sample/ra
      -- 
    ra_927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_190_inst_ack_0, ack => maxPool4_CP_307_elements(114)); -- 
    -- CP-element group 115:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	376 
    -- CP-element group 115: marked-successors 
    -- CP-element group 115: 	113 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 assign_stmt_89_to_assign_stmt_1130/slice_190_update_completed_
      -- CP-element group 115: 	 assign_stmt_89_to_assign_stmt_1130/slice_190_Update/$exit
      -- CP-element group 115: 	 assign_stmt_89_to_assign_stmt_1130/slice_190_Update/ca
      -- 
    ca_932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_190_inst_ack_1, ack => maxPool4_CP_307_elements(115)); -- 
    -- CP-element group 116:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	43 
    -- CP-element group 116: marked-predecessors 
    -- CP-element group 116: 	118 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 assign_stmt_89_to_assign_stmt_1130/slice_194_sample_start_
      -- CP-element group 116: 	 assign_stmt_89_to_assign_stmt_1130/slice_194_Sample/$entry
      -- CP-element group 116: 	 assign_stmt_89_to_assign_stmt_1130/slice_194_Sample/rr
      -- 
    rr_940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(116), ack => slice_194_inst_req_0); -- 
    maxPool4_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(43) & maxPool4_CP_307_elements(118);
      gj_maxPool4_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: marked-predecessors 
    -- CP-element group 117: 	119 
    -- CP-element group 117: 	321 
    -- CP-element group 117: 	386 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	119 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 assign_stmt_89_to_assign_stmt_1130/slice_194_update_start_
      -- CP-element group 117: 	 assign_stmt_89_to_assign_stmt_1130/slice_194_Update/$entry
      -- CP-element group 117: 	 assign_stmt_89_to_assign_stmt_1130/slice_194_Update/cr
      -- 
    cr_945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(117), ack => slice_194_inst_req_1); -- 
    maxPool4_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(119) & maxPool4_CP_307_elements(321) & maxPool4_CP_307_elements(386);
      gj_maxPool4_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: successors 
    -- CP-element group 118: marked-successors 
    -- CP-element group 118: 	41 
    -- CP-element group 118: 	116 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 assign_stmt_89_to_assign_stmt_1130/slice_194_sample_completed_
      -- CP-element group 118: 	 assign_stmt_89_to_assign_stmt_1130/slice_194_Sample/$exit
      -- CP-element group 118: 	 assign_stmt_89_to_assign_stmt_1130/slice_194_Sample/ra
      -- 
    ra_941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_194_inst_ack_0, ack => maxPool4_CP_307_elements(118)); -- 
    -- CP-element group 119:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	117 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	319 
    -- CP-element group 119: 	384 
    -- CP-element group 119: marked-successors 
    -- CP-element group 119: 	117 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 assign_stmt_89_to_assign_stmt_1130/slice_194_update_completed_
      -- CP-element group 119: 	 assign_stmt_89_to_assign_stmt_1130/slice_194_Update/$exit
      -- CP-element group 119: 	 assign_stmt_89_to_assign_stmt_1130/slice_194_Update/ca
      -- 
    ca_946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_194_inst_ack_1, ack => maxPool4_CP_307_elements(119)); -- 
    -- CP-element group 120:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	43 
    -- CP-element group 120: marked-predecessors 
    -- CP-element group 120: 	122 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	122 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 assign_stmt_89_to_assign_stmt_1130/slice_198_sample_start_
      -- CP-element group 120: 	 assign_stmt_89_to_assign_stmt_1130/slice_198_Sample/$entry
      -- CP-element group 120: 	 assign_stmt_89_to_assign_stmt_1130/slice_198_Sample/rr
      -- 
    rr_954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(120), ack => slice_198_inst_req_0); -- 
    maxPool4_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(43) & maxPool4_CP_307_elements(122);
      gj_maxPool4_cp_element_group_120 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: marked-predecessors 
    -- CP-element group 121: 	123 
    -- CP-element group 121: 	321 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	123 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 assign_stmt_89_to_assign_stmt_1130/slice_198_update_start_
      -- CP-element group 121: 	 assign_stmt_89_to_assign_stmt_1130/slice_198_Update/$entry
      -- CP-element group 121: 	 assign_stmt_89_to_assign_stmt_1130/slice_198_Update/cr
      -- 
    cr_959_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_959_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(121), ack => slice_198_inst_req_1); -- 
    maxPool4_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(123) & maxPool4_CP_307_elements(321);
      gj_maxPool4_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	120 
    -- CP-element group 122: successors 
    -- CP-element group 122: marked-successors 
    -- CP-element group 122: 	41 
    -- CP-element group 122: 	120 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 assign_stmt_89_to_assign_stmt_1130/slice_198_sample_completed_
      -- CP-element group 122: 	 assign_stmt_89_to_assign_stmt_1130/slice_198_Sample/$exit
      -- CP-element group 122: 	 assign_stmt_89_to_assign_stmt_1130/slice_198_Sample/ra
      -- 
    ra_955_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_198_inst_ack_0, ack => maxPool4_CP_307_elements(122)); -- 
    -- CP-element group 123:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	121 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	319 
    -- CP-element group 123: marked-successors 
    -- CP-element group 123: 	121 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 assign_stmt_89_to_assign_stmt_1130/slice_198_update_completed_
      -- CP-element group 123: 	 assign_stmt_89_to_assign_stmt_1130/slice_198_Update/$exit
      -- CP-element group 123: 	 assign_stmt_89_to_assign_stmt_1130/slice_198_Update/ca
      -- 
    ca_960_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_198_inst_ack_1, ack => maxPool4_CP_307_elements(123)); -- 
    -- CP-element group 124:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	43 
    -- CP-element group 124: marked-predecessors 
    -- CP-element group 124: 	126 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	126 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 assign_stmt_89_to_assign_stmt_1130/slice_202_sample_start_
      -- CP-element group 124: 	 assign_stmt_89_to_assign_stmt_1130/slice_202_Sample/$entry
      -- CP-element group 124: 	 assign_stmt_89_to_assign_stmt_1130/slice_202_Sample/rr
      -- 
    rr_968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(124), ack => slice_202_inst_req_0); -- 
    maxPool4_cp_element_group_124: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_124"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(43) & maxPool4_CP_307_elements(126);
      gj_maxPool4_cp_element_group_124 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(124), clk => clk, reset => reset); --
    end block;
    -- CP-element group 125:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: marked-predecessors 
    -- CP-element group 125: 	127 
    -- CP-element group 125: 	321 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 assign_stmt_89_to_assign_stmt_1130/slice_202_update_start_
      -- CP-element group 125: 	 assign_stmt_89_to_assign_stmt_1130/slice_202_Update/$entry
      -- CP-element group 125: 	 assign_stmt_89_to_assign_stmt_1130/slice_202_Update/cr
      -- 
    cr_973_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_973_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(125), ack => slice_202_inst_req_1); -- 
    maxPool4_cp_element_group_125: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_125"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(127) & maxPool4_CP_307_elements(321);
      gj_maxPool4_cp_element_group_125 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(125), clk => clk, reset => reset); --
    end block;
    -- CP-element group 126:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	124 
    -- CP-element group 126: successors 
    -- CP-element group 126: marked-successors 
    -- CP-element group 126: 	41 
    -- CP-element group 126: 	124 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 assign_stmt_89_to_assign_stmt_1130/slice_202_sample_completed_
      -- CP-element group 126: 	 assign_stmt_89_to_assign_stmt_1130/slice_202_Sample/$exit
      -- CP-element group 126: 	 assign_stmt_89_to_assign_stmt_1130/slice_202_Sample/ra
      -- 
    ra_969_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_202_inst_ack_0, ack => maxPool4_CP_307_elements(126)); -- 
    -- CP-element group 127:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	125 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	319 
    -- CP-element group 127: marked-successors 
    -- CP-element group 127: 	125 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 assign_stmt_89_to_assign_stmt_1130/slice_202_update_completed_
      -- CP-element group 127: 	 assign_stmt_89_to_assign_stmt_1130/slice_202_Update/$exit
      -- CP-element group 127: 	 assign_stmt_89_to_assign_stmt_1130/slice_202_Update/ca
      -- 
    ca_974_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_202_inst_ack_1, ack => maxPool4_CP_307_elements(127)); -- 
    -- CP-element group 128:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	43 
    -- CP-element group 128: marked-predecessors 
    -- CP-element group 128: 	130 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	130 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 assign_stmt_89_to_assign_stmt_1130/slice_206_sample_start_
      -- CP-element group 128: 	 assign_stmt_89_to_assign_stmt_1130/slice_206_Sample/$entry
      -- CP-element group 128: 	 assign_stmt_89_to_assign_stmt_1130/slice_206_Sample/rr
      -- 
    rr_982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(128), ack => slice_206_inst_req_0); -- 
    maxPool4_cp_element_group_128: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_128"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(43) & maxPool4_CP_307_elements(130);
      gj_maxPool4_cp_element_group_128 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(128), clk => clk, reset => reset); --
    end block;
    -- CP-element group 129:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: marked-predecessors 
    -- CP-element group 129: 	131 
    -- CP-element group 129: 	321 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	131 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 assign_stmt_89_to_assign_stmt_1130/slice_206_update_start_
      -- CP-element group 129: 	 assign_stmt_89_to_assign_stmt_1130/slice_206_Update/$entry
      -- CP-element group 129: 	 assign_stmt_89_to_assign_stmt_1130/slice_206_Update/cr
      -- 
    cr_987_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_987_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(129), ack => slice_206_inst_req_1); -- 
    maxPool4_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(131) & maxPool4_CP_307_elements(321);
      gj_maxPool4_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	128 
    -- CP-element group 130: successors 
    -- CP-element group 130: marked-successors 
    -- CP-element group 130: 	41 
    -- CP-element group 130: 	128 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 assign_stmt_89_to_assign_stmt_1130/slice_206_sample_completed_
      -- CP-element group 130: 	 assign_stmt_89_to_assign_stmt_1130/slice_206_Sample/$exit
      -- CP-element group 130: 	 assign_stmt_89_to_assign_stmt_1130/slice_206_Sample/ra
      -- 
    ra_983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_206_inst_ack_0, ack => maxPool4_CP_307_elements(130)); -- 
    -- CP-element group 131:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	129 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	319 
    -- CP-element group 131: marked-successors 
    -- CP-element group 131: 	129 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 assign_stmt_89_to_assign_stmt_1130/slice_206_update_completed_
      -- CP-element group 131: 	 assign_stmt_89_to_assign_stmt_1130/slice_206_Update/$exit
      -- CP-element group 131: 	 assign_stmt_89_to_assign_stmt_1130/slice_206_Update/ca
      -- 
    ca_988_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_206_inst_ack_1, ack => maxPool4_CP_307_elements(131)); -- 
    -- CP-element group 132:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	43 
    -- CP-element group 132: marked-predecessors 
    -- CP-element group 132: 	134 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 assign_stmt_89_to_assign_stmt_1130/slice_210_Sample/rr
      -- CP-element group 132: 	 assign_stmt_89_to_assign_stmt_1130/slice_210_Sample/$entry
      -- CP-element group 132: 	 assign_stmt_89_to_assign_stmt_1130/slice_210_sample_start_
      -- 
    rr_996_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_996_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(132), ack => slice_210_inst_req_0); -- 
    maxPool4_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(43) & maxPool4_CP_307_elements(134);
      gj_maxPool4_cp_element_group_132 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: marked-predecessors 
    -- CP-element group 133: 	135 
    -- CP-element group 133: 	340 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	135 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 assign_stmt_89_to_assign_stmt_1130/slice_210_Update/cr
      -- CP-element group 133: 	 assign_stmt_89_to_assign_stmt_1130/slice_210_Update/$entry
      -- CP-element group 133: 	 assign_stmt_89_to_assign_stmt_1130/slice_210_update_start_
      -- 
    cr_1001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(133), ack => slice_210_inst_req_1); -- 
    maxPool4_cp_element_group_133: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_133"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(135) & maxPool4_CP_307_elements(340);
      gj_maxPool4_cp_element_group_133 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(133), clk => clk, reset => reset); --
    end block;
    -- CP-element group 134:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134: marked-successors 
    -- CP-element group 134: 	41 
    -- CP-element group 134: 	132 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 assign_stmt_89_to_assign_stmt_1130/slice_210_Sample/ra
      -- CP-element group 134: 	 assign_stmt_89_to_assign_stmt_1130/slice_210_Sample/$exit
      -- CP-element group 134: 	 assign_stmt_89_to_assign_stmt_1130/slice_210_sample_completed_
      -- 
    ra_997_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_210_inst_ack_0, ack => maxPool4_CP_307_elements(134)); -- 
    -- CP-element group 135:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	133 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	338 
    -- CP-element group 135: marked-successors 
    -- CP-element group 135: 	133 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 assign_stmt_89_to_assign_stmt_1130/slice_210_Update/ca
      -- CP-element group 135: 	 assign_stmt_89_to_assign_stmt_1130/slice_210_Update/$exit
      -- CP-element group 135: 	 assign_stmt_89_to_assign_stmt_1130/slice_210_update_completed_
      -- 
    ca_1002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_210_inst_ack_1, ack => maxPool4_CP_307_elements(135)); -- 
    -- CP-element group 136:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	43 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	138 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	138 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 assign_stmt_89_to_assign_stmt_1130/slice_214_Sample/rr
      -- CP-element group 136: 	 assign_stmt_89_to_assign_stmt_1130/slice_214_Sample/$entry
      -- CP-element group 136: 	 assign_stmt_89_to_assign_stmt_1130/slice_214_sample_start_
      -- 
    rr_1010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(136), ack => slice_214_inst_req_0); -- 
    maxPool4_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(43) & maxPool4_CP_307_elements(138);
      gj_maxPool4_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: marked-predecessors 
    -- CP-element group 137: 	139 
    -- CP-element group 137: 	340 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	139 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 assign_stmt_89_to_assign_stmt_1130/slice_214_Update/cr
      -- CP-element group 137: 	 assign_stmt_89_to_assign_stmt_1130/slice_214_Update/$entry
      -- CP-element group 137: 	 assign_stmt_89_to_assign_stmt_1130/slice_214_update_start_
      -- 
    cr_1015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(137), ack => slice_214_inst_req_1); -- 
    maxPool4_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(139) & maxPool4_CP_307_elements(340);
      gj_maxPool4_cp_element_group_137 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	136 
    -- CP-element group 138: successors 
    -- CP-element group 138: marked-successors 
    -- CP-element group 138: 	41 
    -- CP-element group 138: 	136 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 assign_stmt_89_to_assign_stmt_1130/slice_214_Sample/ra
      -- CP-element group 138: 	 assign_stmt_89_to_assign_stmt_1130/slice_214_Sample/$exit
      -- CP-element group 138: 	 assign_stmt_89_to_assign_stmt_1130/slice_214_sample_completed_
      -- 
    ra_1011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_214_inst_ack_0, ack => maxPool4_CP_307_elements(138)); -- 
    -- CP-element group 139:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	137 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	338 
    -- CP-element group 139: marked-successors 
    -- CP-element group 139: 	137 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 assign_stmt_89_to_assign_stmt_1130/slice_214_Update/ca
      -- CP-element group 139: 	 assign_stmt_89_to_assign_stmt_1130/slice_214_Update/$exit
      -- CP-element group 139: 	 assign_stmt_89_to_assign_stmt_1130/slice_214_update_completed_
      -- 
    ca_1016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_214_inst_ack_1, ack => maxPool4_CP_307_elements(139)); -- 
    -- CP-element group 140:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	43 
    -- CP-element group 140: marked-predecessors 
    -- CP-element group 140: 	142 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	142 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 assign_stmt_89_to_assign_stmt_1130/slice_218_sample_start_
      -- CP-element group 140: 	 assign_stmt_89_to_assign_stmt_1130/slice_218_Sample/rr
      -- CP-element group 140: 	 assign_stmt_89_to_assign_stmt_1130/slice_218_Sample/$entry
      -- 
    rr_1024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(140), ack => slice_218_inst_req_0); -- 
    maxPool4_cp_element_group_140: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_140"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(43) & maxPool4_CP_307_elements(142);
      gj_maxPool4_cp_element_group_140 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(140), clk => clk, reset => reset); --
    end block;
    -- CP-element group 141:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: marked-predecessors 
    -- CP-element group 141: 	143 
    -- CP-element group 141: 	340 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	143 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 assign_stmt_89_to_assign_stmt_1130/slice_218_Update/cr
      -- CP-element group 141: 	 assign_stmt_89_to_assign_stmt_1130/slice_218_Update/$entry
      -- CP-element group 141: 	 assign_stmt_89_to_assign_stmt_1130/slice_218_update_start_
      -- 
    cr_1029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(141), ack => slice_218_inst_req_1); -- 
    maxPool4_cp_element_group_141: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_141"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(143) & maxPool4_CP_307_elements(340);
      gj_maxPool4_cp_element_group_141 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(141), clk => clk, reset => reset); --
    end block;
    -- CP-element group 142:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	140 
    -- CP-element group 142: successors 
    -- CP-element group 142: marked-successors 
    -- CP-element group 142: 	41 
    -- CP-element group 142: 	140 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 assign_stmt_89_to_assign_stmt_1130/slice_218_Sample/ra
      -- CP-element group 142: 	 assign_stmt_89_to_assign_stmt_1130/slice_218_Sample/$exit
      -- CP-element group 142: 	 assign_stmt_89_to_assign_stmt_1130/slice_218_sample_completed_
      -- 
    ra_1025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_218_inst_ack_0, ack => maxPool4_CP_307_elements(142)); -- 
    -- CP-element group 143:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	141 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	338 
    -- CP-element group 143: marked-successors 
    -- CP-element group 143: 	141 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 assign_stmt_89_to_assign_stmt_1130/slice_218_Update/ca
      -- CP-element group 143: 	 assign_stmt_89_to_assign_stmt_1130/slice_218_Update/$exit
      -- CP-element group 143: 	 assign_stmt_89_to_assign_stmt_1130/slice_218_update_completed_
      -- 
    ca_1030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_218_inst_ack_1, ack => maxPool4_CP_307_elements(143)); -- 
    -- CP-element group 144:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	43 
    -- CP-element group 144: marked-predecessors 
    -- CP-element group 144: 	146 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	146 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 assign_stmt_89_to_assign_stmt_1130/slice_222_Sample/rr
      -- CP-element group 144: 	 assign_stmt_89_to_assign_stmt_1130/slice_222_Sample/$entry
      -- CP-element group 144: 	 assign_stmt_89_to_assign_stmt_1130/slice_222_sample_start_
      -- 
    rr_1038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(144), ack => slice_222_inst_req_0); -- 
    maxPool4_cp_element_group_144: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_144"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(43) & maxPool4_CP_307_elements(146);
      gj_maxPool4_cp_element_group_144 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(144), clk => clk, reset => reset); --
    end block;
    -- CP-element group 145:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: marked-predecessors 
    -- CP-element group 145: 	147 
    -- CP-element group 145: 	340 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	147 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 assign_stmt_89_to_assign_stmt_1130/slice_222_Update/cr
      -- CP-element group 145: 	 assign_stmt_89_to_assign_stmt_1130/slice_222_Update/$entry
      -- CP-element group 145: 	 assign_stmt_89_to_assign_stmt_1130/slice_222_update_start_
      -- 
    cr_1043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(145), ack => slice_222_inst_req_1); -- 
    maxPool4_cp_element_group_145: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_145"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(147) & maxPool4_CP_307_elements(340);
      gj_maxPool4_cp_element_group_145 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(145), clk => clk, reset => reset); --
    end block;
    -- CP-element group 146:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	144 
    -- CP-element group 146: successors 
    -- CP-element group 146: marked-successors 
    -- CP-element group 146: 	41 
    -- CP-element group 146: 	144 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 assign_stmt_89_to_assign_stmt_1130/slice_222_Sample/ra
      -- CP-element group 146: 	 assign_stmt_89_to_assign_stmt_1130/slice_222_Sample/$exit
      -- CP-element group 146: 	 assign_stmt_89_to_assign_stmt_1130/slice_222_sample_completed_
      -- 
    ra_1039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_222_inst_ack_0, ack => maxPool4_CP_307_elements(146)); -- 
    -- CP-element group 147:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	145 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	338 
    -- CP-element group 147: marked-successors 
    -- CP-element group 147: 	145 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 assign_stmt_89_to_assign_stmt_1130/slice_222_Update/ca
      -- CP-element group 147: 	 assign_stmt_89_to_assign_stmt_1130/slice_222_Update/$exit
      -- CP-element group 147: 	 assign_stmt_89_to_assign_stmt_1130/slice_222_update_completed_
      -- 
    ca_1044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_222_inst_ack_1, ack => maxPool4_CP_307_elements(147)); -- 
    -- CP-element group 148:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	43 
    -- CP-element group 148: marked-predecessors 
    -- CP-element group 148: 	150 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	150 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 assign_stmt_89_to_assign_stmt_1130/slice_226_Sample/rr
      -- CP-element group 148: 	 assign_stmt_89_to_assign_stmt_1130/slice_226_Sample/$entry
      -- CP-element group 148: 	 assign_stmt_89_to_assign_stmt_1130/slice_226_sample_start_
      -- 
    rr_1052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(148), ack => slice_226_inst_req_0); -- 
    maxPool4_cp_element_group_148: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_148"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(43) & maxPool4_CP_307_elements(150);
      gj_maxPool4_cp_element_group_148 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(148), clk => clk, reset => reset); --
    end block;
    -- CP-element group 149:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: marked-predecessors 
    -- CP-element group 149: 	151 
    -- CP-element group 149: 	359 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	151 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 assign_stmt_89_to_assign_stmt_1130/slice_226_Update/$entry
      -- CP-element group 149: 	 assign_stmt_89_to_assign_stmt_1130/slice_226_update_start_
      -- CP-element group 149: 	 assign_stmt_89_to_assign_stmt_1130/slice_226_Update/cr
      -- 
    cr_1057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(149), ack => slice_226_inst_req_1); -- 
    maxPool4_cp_element_group_149: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_149"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(151) & maxPool4_CP_307_elements(359);
      gj_maxPool4_cp_element_group_149 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(149), clk => clk, reset => reset); --
    end block;
    -- CP-element group 150:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	148 
    -- CP-element group 150: successors 
    -- CP-element group 150: marked-successors 
    -- CP-element group 150: 	41 
    -- CP-element group 150: 	148 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 assign_stmt_89_to_assign_stmt_1130/slice_226_Sample/ra
      -- CP-element group 150: 	 assign_stmt_89_to_assign_stmt_1130/slice_226_Sample/$exit
      -- CP-element group 150: 	 assign_stmt_89_to_assign_stmt_1130/slice_226_sample_completed_
      -- 
    ra_1053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_226_inst_ack_0, ack => maxPool4_CP_307_elements(150)); -- 
    -- CP-element group 151:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	149 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	357 
    -- CP-element group 151: marked-successors 
    -- CP-element group 151: 	149 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 assign_stmt_89_to_assign_stmt_1130/slice_226_Update/$exit
      -- CP-element group 151: 	 assign_stmt_89_to_assign_stmt_1130/slice_226_update_completed_
      -- CP-element group 151: 	 assign_stmt_89_to_assign_stmt_1130/slice_226_Update/ca
      -- 
    ca_1058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_226_inst_ack_1, ack => maxPool4_CP_307_elements(151)); -- 
    -- CP-element group 152:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	43 
    -- CP-element group 152: marked-predecessors 
    -- CP-element group 152: 	154 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	154 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 assign_stmt_89_to_assign_stmt_1130/slice_230_Sample/rr
      -- CP-element group 152: 	 assign_stmt_89_to_assign_stmt_1130/slice_230_Sample/$entry
      -- CP-element group 152: 	 assign_stmt_89_to_assign_stmt_1130/slice_230_sample_start_
      -- 
    rr_1066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(152), ack => slice_230_inst_req_0); -- 
    maxPool4_cp_element_group_152: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_152"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(43) & maxPool4_CP_307_elements(154);
      gj_maxPool4_cp_element_group_152 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(152), clk => clk, reset => reset); --
    end block;
    -- CP-element group 153:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: marked-predecessors 
    -- CP-element group 153: 	155 
    -- CP-element group 153: 	359 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	155 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 assign_stmt_89_to_assign_stmt_1130/slice_230_Update/cr
      -- CP-element group 153: 	 assign_stmt_89_to_assign_stmt_1130/slice_230_Update/$entry
      -- CP-element group 153: 	 assign_stmt_89_to_assign_stmt_1130/slice_230_update_start_
      -- 
    cr_1071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(153), ack => slice_230_inst_req_1); -- 
    maxPool4_cp_element_group_153: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_153"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(155) & maxPool4_CP_307_elements(359);
      gj_maxPool4_cp_element_group_153 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(153), clk => clk, reset => reset); --
    end block;
    -- CP-element group 154:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	152 
    -- CP-element group 154: successors 
    -- CP-element group 154: marked-successors 
    -- CP-element group 154: 	41 
    -- CP-element group 154: 	152 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 assign_stmt_89_to_assign_stmt_1130/slice_230_Sample/ra
      -- CP-element group 154: 	 assign_stmt_89_to_assign_stmt_1130/slice_230_Sample/$exit
      -- CP-element group 154: 	 assign_stmt_89_to_assign_stmt_1130/slice_230_sample_completed_
      -- 
    ra_1067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_230_inst_ack_0, ack => maxPool4_CP_307_elements(154)); -- 
    -- CP-element group 155:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	153 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	357 
    -- CP-element group 155: marked-successors 
    -- CP-element group 155: 	153 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 assign_stmt_89_to_assign_stmt_1130/slice_230_Update/ca
      -- CP-element group 155: 	 assign_stmt_89_to_assign_stmt_1130/slice_230_Update/$exit
      -- CP-element group 155: 	 assign_stmt_89_to_assign_stmt_1130/slice_230_update_completed_
      -- 
    ca_1072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_230_inst_ack_1, ack => maxPool4_CP_307_elements(155)); -- 
    -- CP-element group 156:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	43 
    -- CP-element group 156: marked-predecessors 
    -- CP-element group 156: 	158 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 assign_stmt_89_to_assign_stmt_1130/slice_234_Sample/rr
      -- CP-element group 156: 	 assign_stmt_89_to_assign_stmt_1130/slice_234_Sample/$entry
      -- CP-element group 156: 	 assign_stmt_89_to_assign_stmt_1130/slice_234_sample_start_
      -- 
    rr_1080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(156), ack => slice_234_inst_req_0); -- 
    maxPool4_cp_element_group_156: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_156"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(43) & maxPool4_CP_307_elements(158);
      gj_maxPool4_cp_element_group_156 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(156), clk => clk, reset => reset); --
    end block;
    -- CP-element group 157:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: marked-predecessors 
    -- CP-element group 157: 	159 
    -- CP-element group 157: 	359 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	159 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 assign_stmt_89_to_assign_stmt_1130/slice_234_Update/$entry
      -- CP-element group 157: 	 assign_stmt_89_to_assign_stmt_1130/slice_234_update_start_
      -- CP-element group 157: 	 assign_stmt_89_to_assign_stmt_1130/slice_234_Update/cr
      -- 
    cr_1085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(157), ack => slice_234_inst_req_1); -- 
    maxPool4_cp_element_group_157: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_157"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(159) & maxPool4_CP_307_elements(359);
      gj_maxPool4_cp_element_group_157 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(157), clk => clk, reset => reset); --
    end block;
    -- CP-element group 158:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	156 
    -- CP-element group 158: successors 
    -- CP-element group 158: marked-successors 
    -- CP-element group 158: 	41 
    -- CP-element group 158: 	156 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 assign_stmt_89_to_assign_stmt_1130/slice_234_Sample/ra
      -- CP-element group 158: 	 assign_stmt_89_to_assign_stmt_1130/slice_234_Sample/$exit
      -- CP-element group 158: 	 assign_stmt_89_to_assign_stmt_1130/slice_234_sample_completed_
      -- 
    ra_1081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_234_inst_ack_0, ack => maxPool4_CP_307_elements(158)); -- 
    -- CP-element group 159:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	157 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	357 
    -- CP-element group 159: marked-successors 
    -- CP-element group 159: 	157 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 assign_stmt_89_to_assign_stmt_1130/slice_234_update_completed_
      -- CP-element group 159: 	 assign_stmt_89_to_assign_stmt_1130/slice_234_Update/ca
      -- CP-element group 159: 	 assign_stmt_89_to_assign_stmt_1130/slice_234_Update/$exit
      -- 
    ca_1086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_234_inst_ack_1, ack => maxPool4_CP_307_elements(159)); -- 
    -- CP-element group 160:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	43 
    -- CP-element group 160: marked-predecessors 
    -- CP-element group 160: 	162 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	162 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 assign_stmt_89_to_assign_stmt_1130/slice_238_Sample/rr
      -- CP-element group 160: 	 assign_stmt_89_to_assign_stmt_1130/slice_238_Sample/$entry
      -- CP-element group 160: 	 assign_stmt_89_to_assign_stmt_1130/slice_238_sample_start_
      -- 
    rr_1094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(160), ack => slice_238_inst_req_0); -- 
    maxPool4_cp_element_group_160: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_160"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(43) & maxPool4_CP_307_elements(162);
      gj_maxPool4_cp_element_group_160 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(160), clk => clk, reset => reset); --
    end block;
    -- CP-element group 161:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: marked-predecessors 
    -- CP-element group 161: 	163 
    -- CP-element group 161: 	359 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	163 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 assign_stmt_89_to_assign_stmt_1130/slice_238_Update/cr
      -- CP-element group 161: 	 assign_stmt_89_to_assign_stmt_1130/slice_238_Update/$entry
      -- CP-element group 161: 	 assign_stmt_89_to_assign_stmt_1130/slice_238_update_start_
      -- 
    cr_1099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(161), ack => slice_238_inst_req_1); -- 
    maxPool4_cp_element_group_161: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_161"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(163) & maxPool4_CP_307_elements(359);
      gj_maxPool4_cp_element_group_161 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(161), clk => clk, reset => reset); --
    end block;
    -- CP-element group 162:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	160 
    -- CP-element group 162: successors 
    -- CP-element group 162: marked-successors 
    -- CP-element group 162: 	41 
    -- CP-element group 162: 	160 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 assign_stmt_89_to_assign_stmt_1130/slice_238_Sample/ra
      -- CP-element group 162: 	 assign_stmt_89_to_assign_stmt_1130/slice_238_Sample/$exit
      -- CP-element group 162: 	 assign_stmt_89_to_assign_stmt_1130/slice_238_sample_completed_
      -- 
    ra_1095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_238_inst_ack_0, ack => maxPool4_CP_307_elements(162)); -- 
    -- CP-element group 163:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	161 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	357 
    -- CP-element group 163: marked-successors 
    -- CP-element group 163: 	161 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 assign_stmt_89_to_assign_stmt_1130/slice_238_Update/ca
      -- CP-element group 163: 	 assign_stmt_89_to_assign_stmt_1130/slice_238_Update/$exit
      -- CP-element group 163: 	 assign_stmt_89_to_assign_stmt_1130/slice_238_update_completed_
      -- 
    ca_1100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_238_inst_ack_1, ack => maxPool4_CP_307_elements(163)); -- 
    -- CP-element group 164:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	43 
    -- CP-element group 164: marked-predecessors 
    -- CP-element group 164: 	166 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 assign_stmt_89_to_assign_stmt_1130/slice_242_Sample/$entry
      -- CP-element group 164: 	 assign_stmt_89_to_assign_stmt_1130/slice_242_Sample/rr
      -- CP-element group 164: 	 assign_stmt_89_to_assign_stmt_1130/slice_242_sample_start_
      -- 
    rr_1108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(164), ack => slice_242_inst_req_0); -- 
    maxPool4_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(43) & maxPool4_CP_307_elements(166);
      gj_maxPool4_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: marked-predecessors 
    -- CP-element group 165: 	167 
    -- CP-element group 165: 	378 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	167 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 assign_stmt_89_to_assign_stmt_1130/slice_242_Update/cr
      -- CP-element group 165: 	 assign_stmt_89_to_assign_stmt_1130/slice_242_update_start_
      -- CP-element group 165: 	 assign_stmt_89_to_assign_stmt_1130/slice_242_Update/$entry
      -- 
    cr_1113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(165), ack => slice_242_inst_req_1); -- 
    maxPool4_cp_element_group_165: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_165"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(167) & maxPool4_CP_307_elements(378);
      gj_maxPool4_cp_element_group_165 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(165), clk => clk, reset => reset); --
    end block;
    -- CP-element group 166:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: successors 
    -- CP-element group 166: marked-successors 
    -- CP-element group 166: 	41 
    -- CP-element group 166: 	164 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 assign_stmt_89_to_assign_stmt_1130/slice_242_Sample/$exit
      -- CP-element group 166: 	 assign_stmt_89_to_assign_stmt_1130/slice_242_sample_completed_
      -- CP-element group 166: 	 assign_stmt_89_to_assign_stmt_1130/slice_242_Sample/ra
      -- 
    ra_1109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_242_inst_ack_0, ack => maxPool4_CP_307_elements(166)); -- 
    -- CP-element group 167:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	165 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	376 
    -- CP-element group 167: marked-successors 
    -- CP-element group 167: 	165 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 assign_stmt_89_to_assign_stmt_1130/slice_242_update_completed_
      -- CP-element group 167: 	 assign_stmt_89_to_assign_stmt_1130/slice_242_Update/$exit
      -- CP-element group 167: 	 assign_stmt_89_to_assign_stmt_1130/slice_242_Update/ca
      -- 
    ca_1114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_242_inst_ack_1, ack => maxPool4_CP_307_elements(167)); -- 
    -- CP-element group 168:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	43 
    -- CP-element group 168: marked-predecessors 
    -- CP-element group 168: 	170 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	170 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 assign_stmt_89_to_assign_stmt_1130/slice_246_sample_start_
      -- CP-element group 168: 	 assign_stmt_89_to_assign_stmt_1130/slice_246_Sample/rr
      -- CP-element group 168: 	 assign_stmt_89_to_assign_stmt_1130/slice_246_Sample/$entry
      -- 
    rr_1122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(168), ack => slice_246_inst_req_0); -- 
    maxPool4_cp_element_group_168: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_168"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(43) & maxPool4_CP_307_elements(170);
      gj_maxPool4_cp_element_group_168 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(168), clk => clk, reset => reset); --
    end block;
    -- CP-element group 169:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: marked-predecessors 
    -- CP-element group 169: 	171 
    -- CP-element group 169: 	378 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	171 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 assign_stmt_89_to_assign_stmt_1130/slice_246_Update/$entry
      -- CP-element group 169: 	 assign_stmt_89_to_assign_stmt_1130/slice_246_update_start_
      -- CP-element group 169: 	 assign_stmt_89_to_assign_stmt_1130/slice_246_Update/cr
      -- 
    cr_1127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(169), ack => slice_246_inst_req_1); -- 
    maxPool4_cp_element_group_169: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_169"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(171) & maxPool4_CP_307_elements(378);
      gj_maxPool4_cp_element_group_169 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(169), clk => clk, reset => reset); --
    end block;
    -- CP-element group 170:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	168 
    -- CP-element group 170: successors 
    -- CP-element group 170: marked-successors 
    -- CP-element group 170: 	41 
    -- CP-element group 170: 	168 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 assign_stmt_89_to_assign_stmt_1130/slice_246_Sample/ra
      -- CP-element group 170: 	 assign_stmt_89_to_assign_stmt_1130/slice_246_Sample/$exit
      -- CP-element group 170: 	 assign_stmt_89_to_assign_stmt_1130/slice_246_sample_completed_
      -- 
    ra_1123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_246_inst_ack_0, ack => maxPool4_CP_307_elements(170)); -- 
    -- CP-element group 171:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	169 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	376 
    -- CP-element group 171: marked-successors 
    -- CP-element group 171: 	169 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 assign_stmt_89_to_assign_stmt_1130/slice_246_Update/$exit
      -- CP-element group 171: 	 assign_stmt_89_to_assign_stmt_1130/slice_246_update_completed_
      -- CP-element group 171: 	 assign_stmt_89_to_assign_stmt_1130/slice_246_Update/ca
      -- 
    ca_1128_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_246_inst_ack_1, ack => maxPool4_CP_307_elements(171)); -- 
    -- CP-element group 172:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	43 
    -- CP-element group 172: marked-predecessors 
    -- CP-element group 172: 	174 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	174 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 assign_stmt_89_to_assign_stmt_1130/slice_250_Sample/$entry
      -- CP-element group 172: 	 assign_stmt_89_to_assign_stmt_1130/slice_250_sample_start_
      -- CP-element group 172: 	 assign_stmt_89_to_assign_stmt_1130/slice_250_Sample/rr
      -- 
    rr_1136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(172), ack => slice_250_inst_req_0); -- 
    maxPool4_cp_element_group_172: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_172"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(43) & maxPool4_CP_307_elements(174);
      gj_maxPool4_cp_element_group_172 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(172), clk => clk, reset => reset); --
    end block;
    -- CP-element group 173:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: marked-predecessors 
    -- CP-element group 173: 	175 
    -- CP-element group 173: 	378 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	175 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 assign_stmt_89_to_assign_stmt_1130/slice_250_update_start_
      -- CP-element group 173: 	 assign_stmt_89_to_assign_stmt_1130/slice_250_Update/$entry
      -- CP-element group 173: 	 assign_stmt_89_to_assign_stmt_1130/slice_250_Update/cr
      -- 
    cr_1141_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1141_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(173), ack => slice_250_inst_req_1); -- 
    maxPool4_cp_element_group_173: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_173"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(175) & maxPool4_CP_307_elements(378);
      gj_maxPool4_cp_element_group_173 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(173), clk => clk, reset => reset); --
    end block;
    -- CP-element group 174:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	172 
    -- CP-element group 174: successors 
    -- CP-element group 174: marked-successors 
    -- CP-element group 174: 	41 
    -- CP-element group 174: 	172 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 assign_stmt_89_to_assign_stmt_1130/slice_250_Sample/$exit
      -- CP-element group 174: 	 assign_stmt_89_to_assign_stmt_1130/slice_250_sample_completed_
      -- CP-element group 174: 	 assign_stmt_89_to_assign_stmt_1130/slice_250_Sample/ra
      -- 
    ra_1137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_250_inst_ack_0, ack => maxPool4_CP_307_elements(174)); -- 
    -- CP-element group 175:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	173 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	376 
    -- CP-element group 175: marked-successors 
    -- CP-element group 175: 	173 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 assign_stmt_89_to_assign_stmt_1130/slice_250_update_completed_
      -- CP-element group 175: 	 assign_stmt_89_to_assign_stmt_1130/slice_250_Update/$exit
      -- CP-element group 175: 	 assign_stmt_89_to_assign_stmt_1130/slice_250_Update/ca
      -- 
    ca_1142_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_250_inst_ack_1, ack => maxPool4_CP_307_elements(175)); -- 
    -- CP-element group 176:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	43 
    -- CP-element group 176: marked-predecessors 
    -- CP-element group 176: 	178 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	178 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 assign_stmt_89_to_assign_stmt_1130/slice_254_sample_start_
      -- CP-element group 176: 	 assign_stmt_89_to_assign_stmt_1130/slice_254_Sample/rr
      -- CP-element group 176: 	 assign_stmt_89_to_assign_stmt_1130/slice_254_Sample/$entry
      -- 
    rr_1150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(176), ack => slice_254_inst_req_0); -- 
    maxPool4_cp_element_group_176: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_176"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(43) & maxPool4_CP_307_elements(178);
      gj_maxPool4_cp_element_group_176 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(176), clk => clk, reset => reset); --
    end block;
    -- CP-element group 177:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: marked-predecessors 
    -- CP-element group 177: 	179 
    -- CP-element group 177: 	378 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	179 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 assign_stmt_89_to_assign_stmt_1130/slice_254_Update/cr
      -- CP-element group 177: 	 assign_stmt_89_to_assign_stmt_1130/slice_254_Update/$entry
      -- CP-element group 177: 	 assign_stmt_89_to_assign_stmt_1130/slice_254_update_start_
      -- 
    cr_1155_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1155_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(177), ack => slice_254_inst_req_1); -- 
    maxPool4_cp_element_group_177: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_177"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(179) & maxPool4_CP_307_elements(378);
      gj_maxPool4_cp_element_group_177 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(177), clk => clk, reset => reset); --
    end block;
    -- CP-element group 178:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	176 
    -- CP-element group 178: successors 
    -- CP-element group 178: marked-successors 
    -- CP-element group 178: 	41 
    -- CP-element group 178: 	176 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 assign_stmt_89_to_assign_stmt_1130/slice_254_sample_completed_
      -- CP-element group 178: 	 assign_stmt_89_to_assign_stmt_1130/slice_254_Sample/ra
      -- CP-element group 178: 	 assign_stmt_89_to_assign_stmt_1130/slice_254_Sample/$exit
      -- 
    ra_1151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_254_inst_ack_0, ack => maxPool4_CP_307_elements(178)); -- 
    -- CP-element group 179:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	177 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	376 
    -- CP-element group 179: marked-successors 
    -- CP-element group 179: 	177 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 assign_stmt_89_to_assign_stmt_1130/slice_254_Update/ca
      -- CP-element group 179: 	 assign_stmt_89_to_assign_stmt_1130/slice_254_Update/$exit
      -- CP-element group 179: 	 assign_stmt_89_to_assign_stmt_1130/slice_254_update_completed_
      -- 
    ca_1156_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_254_inst_ack_1, ack => maxPool4_CP_307_elements(179)); -- 
    -- CP-element group 180:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	47 
    -- CP-element group 180: marked-predecessors 
    -- CP-element group 180: 	182 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	182 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 assign_stmt_89_to_assign_stmt_1130/slice_258_sample_start_
      -- CP-element group 180: 	 assign_stmt_89_to_assign_stmt_1130/slice_258_Sample/$entry
      -- CP-element group 180: 	 assign_stmt_89_to_assign_stmt_1130/slice_258_Sample/rr
      -- 
    rr_1164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(180), ack => slice_258_inst_req_0); -- 
    maxPool4_cp_element_group_180: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_180"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(47) & maxPool4_CP_307_elements(182);
      gj_maxPool4_cp_element_group_180 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(180), clk => clk, reset => reset); --
    end block;
    -- CP-element group 181:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: marked-predecessors 
    -- CP-element group 181: 	183 
    -- CP-element group 181: 	321 
    -- CP-element group 181: 	386 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	183 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 assign_stmt_89_to_assign_stmt_1130/slice_258_Update/cr
      -- CP-element group 181: 	 assign_stmt_89_to_assign_stmt_1130/slice_258_Update/$entry
      -- CP-element group 181: 	 assign_stmt_89_to_assign_stmt_1130/slice_258_update_start_
      -- 
    cr_1169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(181), ack => slice_258_inst_req_1); -- 
    maxPool4_cp_element_group_181: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_181"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(183) & maxPool4_CP_307_elements(321) & maxPool4_CP_307_elements(386);
      gj_maxPool4_cp_element_group_181 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(181), clk => clk, reset => reset); --
    end block;
    -- CP-element group 182:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	180 
    -- CP-element group 182: successors 
    -- CP-element group 182: marked-successors 
    -- CP-element group 182: 	45 
    -- CP-element group 182: 	180 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 assign_stmt_89_to_assign_stmt_1130/slice_258_sample_completed_
      -- CP-element group 182: 	 assign_stmt_89_to_assign_stmt_1130/slice_258_Sample/ra
      -- CP-element group 182: 	 assign_stmt_89_to_assign_stmt_1130/slice_258_Sample/$exit
      -- 
    ra_1165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_258_inst_ack_0, ack => maxPool4_CP_307_elements(182)); -- 
    -- CP-element group 183:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	181 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	319 
    -- CP-element group 183: 	384 
    -- CP-element group 183: marked-successors 
    -- CP-element group 183: 	181 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 assign_stmt_89_to_assign_stmt_1130/slice_258_update_completed_
      -- CP-element group 183: 	 assign_stmt_89_to_assign_stmt_1130/slice_258_Update/ca
      -- CP-element group 183: 	 assign_stmt_89_to_assign_stmt_1130/slice_258_Update/$exit
      -- 
    ca_1170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_258_inst_ack_1, ack => maxPool4_CP_307_elements(183)); -- 
    -- CP-element group 184:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	47 
    -- CP-element group 184: marked-predecessors 
    -- CP-element group 184: 	186 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	186 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 assign_stmt_89_to_assign_stmt_1130/slice_262_sample_start_
      -- CP-element group 184: 	 assign_stmt_89_to_assign_stmt_1130/slice_262_Sample/rr
      -- CP-element group 184: 	 assign_stmt_89_to_assign_stmt_1130/slice_262_Sample/$entry
      -- 
    rr_1178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(184), ack => slice_262_inst_req_0); -- 
    maxPool4_cp_element_group_184: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_184"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(47) & maxPool4_CP_307_elements(186);
      gj_maxPool4_cp_element_group_184 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(184), clk => clk, reset => reset); --
    end block;
    -- CP-element group 185:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: marked-predecessors 
    -- CP-element group 185: 	187 
    -- CP-element group 185: 	321 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	187 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 assign_stmt_89_to_assign_stmt_1130/slice_262_update_start_
      -- CP-element group 185: 	 assign_stmt_89_to_assign_stmt_1130/slice_262_Update/cr
      -- CP-element group 185: 	 assign_stmt_89_to_assign_stmt_1130/slice_262_Update/$entry
      -- 
    cr_1183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(185), ack => slice_262_inst_req_1); -- 
    maxPool4_cp_element_group_185: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_185"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(187) & maxPool4_CP_307_elements(321);
      gj_maxPool4_cp_element_group_185 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(185), clk => clk, reset => reset); --
    end block;
    -- CP-element group 186:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	184 
    -- CP-element group 186: successors 
    -- CP-element group 186: marked-successors 
    -- CP-element group 186: 	45 
    -- CP-element group 186: 	184 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 assign_stmt_89_to_assign_stmt_1130/slice_262_sample_completed_
      -- CP-element group 186: 	 assign_stmt_89_to_assign_stmt_1130/slice_262_Sample/ra
      -- CP-element group 186: 	 assign_stmt_89_to_assign_stmt_1130/slice_262_Sample/$exit
      -- 
    ra_1179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_262_inst_ack_0, ack => maxPool4_CP_307_elements(186)); -- 
    -- CP-element group 187:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	185 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	319 
    -- CP-element group 187: marked-successors 
    -- CP-element group 187: 	185 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 assign_stmt_89_to_assign_stmt_1130/slice_262_update_completed_
      -- CP-element group 187: 	 assign_stmt_89_to_assign_stmt_1130/slice_262_Update/$exit
      -- CP-element group 187: 	 assign_stmt_89_to_assign_stmt_1130/slice_262_Update/ca
      -- 
    ca_1184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_262_inst_ack_1, ack => maxPool4_CP_307_elements(187)); -- 
    -- CP-element group 188:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	47 
    -- CP-element group 188: marked-predecessors 
    -- CP-element group 188: 	190 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	190 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 assign_stmt_89_to_assign_stmt_1130/slice_266_sample_start_
      -- CP-element group 188: 	 assign_stmt_89_to_assign_stmt_1130/slice_266_Sample/$entry
      -- CP-element group 188: 	 assign_stmt_89_to_assign_stmt_1130/slice_266_Sample/rr
      -- 
    rr_1192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(188), ack => slice_266_inst_req_0); -- 
    maxPool4_cp_element_group_188: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_188"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(47) & maxPool4_CP_307_elements(190);
      gj_maxPool4_cp_element_group_188 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(188), clk => clk, reset => reset); --
    end block;
    -- CP-element group 189:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: marked-predecessors 
    -- CP-element group 189: 	191 
    -- CP-element group 189: 	321 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	191 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 assign_stmt_89_to_assign_stmt_1130/slice_266_update_start_
      -- CP-element group 189: 	 assign_stmt_89_to_assign_stmt_1130/slice_266_Update/cr
      -- CP-element group 189: 	 assign_stmt_89_to_assign_stmt_1130/slice_266_Update/$entry
      -- 
    cr_1197_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1197_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(189), ack => slice_266_inst_req_1); -- 
    maxPool4_cp_element_group_189: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_189"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(191) & maxPool4_CP_307_elements(321);
      gj_maxPool4_cp_element_group_189 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(189), clk => clk, reset => reset); --
    end block;
    -- CP-element group 190:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	188 
    -- CP-element group 190: successors 
    -- CP-element group 190: marked-successors 
    -- CP-element group 190: 	45 
    -- CP-element group 190: 	188 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 assign_stmt_89_to_assign_stmt_1130/slice_266_sample_completed_
      -- CP-element group 190: 	 assign_stmt_89_to_assign_stmt_1130/slice_266_Sample/$exit
      -- CP-element group 190: 	 assign_stmt_89_to_assign_stmt_1130/slice_266_Sample/ra
      -- 
    ra_1193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_266_inst_ack_0, ack => maxPool4_CP_307_elements(190)); -- 
    -- CP-element group 191:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	189 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	319 
    -- CP-element group 191: marked-successors 
    -- CP-element group 191: 	189 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 assign_stmt_89_to_assign_stmt_1130/slice_266_Update/ca
      -- CP-element group 191: 	 assign_stmt_89_to_assign_stmt_1130/slice_266_update_completed_
      -- CP-element group 191: 	 assign_stmt_89_to_assign_stmt_1130/slice_266_Update/$exit
      -- 
    ca_1198_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_266_inst_ack_1, ack => maxPool4_CP_307_elements(191)); -- 
    -- CP-element group 192:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	47 
    -- CP-element group 192: marked-predecessors 
    -- CP-element group 192: 	194 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	194 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 assign_stmt_89_to_assign_stmt_1130/slice_270_Sample/$entry
      -- CP-element group 192: 	 assign_stmt_89_to_assign_stmt_1130/slice_270_Sample/rr
      -- CP-element group 192: 	 assign_stmt_89_to_assign_stmt_1130/slice_270_sample_start_
      -- 
    rr_1206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(192), ack => slice_270_inst_req_0); -- 
    maxPool4_cp_element_group_192: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_192"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(47) & maxPool4_CP_307_elements(194);
      gj_maxPool4_cp_element_group_192 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(192), clk => clk, reset => reset); --
    end block;
    -- CP-element group 193:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: marked-predecessors 
    -- CP-element group 193: 	195 
    -- CP-element group 193: 	321 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	195 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 assign_stmt_89_to_assign_stmt_1130/slice_270_Update/cr
      -- CP-element group 193: 	 assign_stmt_89_to_assign_stmt_1130/slice_270_update_start_
      -- CP-element group 193: 	 assign_stmt_89_to_assign_stmt_1130/slice_270_Update/$entry
      -- 
    cr_1211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(193), ack => slice_270_inst_req_1); -- 
    maxPool4_cp_element_group_193: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_193"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(195) & maxPool4_CP_307_elements(321);
      gj_maxPool4_cp_element_group_193 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(193), clk => clk, reset => reset); --
    end block;
    -- CP-element group 194:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	192 
    -- CP-element group 194: successors 
    -- CP-element group 194: marked-successors 
    -- CP-element group 194: 	45 
    -- CP-element group 194: 	192 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 assign_stmt_89_to_assign_stmt_1130/slice_270_Sample/$exit
      -- CP-element group 194: 	 assign_stmt_89_to_assign_stmt_1130/slice_270_sample_completed_
      -- CP-element group 194: 	 assign_stmt_89_to_assign_stmt_1130/slice_270_Sample/ra
      -- 
    ra_1207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_270_inst_ack_0, ack => maxPool4_CP_307_elements(194)); -- 
    -- CP-element group 195:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	193 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	319 
    -- CP-element group 195: marked-successors 
    -- CP-element group 195: 	193 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 assign_stmt_89_to_assign_stmt_1130/slice_270_Update/ca
      -- CP-element group 195: 	 assign_stmt_89_to_assign_stmt_1130/slice_270_update_completed_
      -- CP-element group 195: 	 assign_stmt_89_to_assign_stmt_1130/slice_270_Update/$exit
      -- 
    ca_1212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_270_inst_ack_1, ack => maxPool4_CP_307_elements(195)); -- 
    -- CP-element group 196:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	47 
    -- CP-element group 196: marked-predecessors 
    -- CP-element group 196: 	198 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	198 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 assign_stmt_89_to_assign_stmt_1130/slice_274_sample_start_
      -- CP-element group 196: 	 assign_stmt_89_to_assign_stmt_1130/slice_274_Sample/$entry
      -- CP-element group 196: 	 assign_stmt_89_to_assign_stmt_1130/slice_274_Sample/rr
      -- 
    rr_1220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(196), ack => slice_274_inst_req_0); -- 
    maxPool4_cp_element_group_196: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_196"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(47) & maxPool4_CP_307_elements(198);
      gj_maxPool4_cp_element_group_196 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(196), clk => clk, reset => reset); --
    end block;
    -- CP-element group 197:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: marked-predecessors 
    -- CP-element group 197: 	199 
    -- CP-element group 197: 	340 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	199 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 assign_stmt_89_to_assign_stmt_1130/slice_274_Update/$entry
      -- CP-element group 197: 	 assign_stmt_89_to_assign_stmt_1130/slice_274_update_start_
      -- CP-element group 197: 	 assign_stmt_89_to_assign_stmt_1130/slice_274_Update/cr
      -- 
    cr_1225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(197), ack => slice_274_inst_req_1); -- 
    maxPool4_cp_element_group_197: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_197"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(199) & maxPool4_CP_307_elements(340);
      gj_maxPool4_cp_element_group_197 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(197), clk => clk, reset => reset); --
    end block;
    -- CP-element group 198:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	196 
    -- CP-element group 198: successors 
    -- CP-element group 198: marked-successors 
    -- CP-element group 198: 	45 
    -- CP-element group 198: 	196 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 assign_stmt_89_to_assign_stmt_1130/slice_274_Sample/ra
      -- CP-element group 198: 	 assign_stmt_89_to_assign_stmt_1130/slice_274_sample_completed_
      -- CP-element group 198: 	 assign_stmt_89_to_assign_stmt_1130/slice_274_Sample/$exit
      -- 
    ra_1221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_274_inst_ack_0, ack => maxPool4_CP_307_elements(198)); -- 
    -- CP-element group 199:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	197 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	338 
    -- CP-element group 199: marked-successors 
    -- CP-element group 199: 	197 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 assign_stmt_89_to_assign_stmt_1130/slice_274_Update/$exit
      -- CP-element group 199: 	 assign_stmt_89_to_assign_stmt_1130/slice_274_update_completed_
      -- CP-element group 199: 	 assign_stmt_89_to_assign_stmt_1130/slice_274_Update/ca
      -- 
    ca_1226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_274_inst_ack_1, ack => maxPool4_CP_307_elements(199)); -- 
    -- CP-element group 200:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	47 
    -- CP-element group 200: marked-predecessors 
    -- CP-element group 200: 	202 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	202 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 assign_stmt_89_to_assign_stmt_1130/slice_278_sample_start_
      -- CP-element group 200: 	 assign_stmt_89_to_assign_stmt_1130/slice_278_Sample/$entry
      -- CP-element group 200: 	 assign_stmt_89_to_assign_stmt_1130/slice_278_Sample/rr
      -- 
    rr_1234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(200), ack => slice_278_inst_req_0); -- 
    maxPool4_cp_element_group_200: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_200"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(47) & maxPool4_CP_307_elements(202);
      gj_maxPool4_cp_element_group_200 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(200), clk => clk, reset => reset); --
    end block;
    -- CP-element group 201:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: marked-predecessors 
    -- CP-element group 201: 	203 
    -- CP-element group 201: 	340 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	203 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 assign_stmt_89_to_assign_stmt_1130/slice_278_update_start_
      -- CP-element group 201: 	 assign_stmt_89_to_assign_stmt_1130/slice_278_Update/$entry
      -- CP-element group 201: 	 assign_stmt_89_to_assign_stmt_1130/slice_278_Update/cr
      -- 
    cr_1239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(201), ack => slice_278_inst_req_1); -- 
    maxPool4_cp_element_group_201: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_201"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(203) & maxPool4_CP_307_elements(340);
      gj_maxPool4_cp_element_group_201 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(201), clk => clk, reset => reset); --
    end block;
    -- CP-element group 202:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	200 
    -- CP-element group 202: successors 
    -- CP-element group 202: marked-successors 
    -- CP-element group 202: 	45 
    -- CP-element group 202: 	200 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 assign_stmt_89_to_assign_stmt_1130/slice_278_sample_completed_
      -- CP-element group 202: 	 assign_stmt_89_to_assign_stmt_1130/slice_278_Sample/$exit
      -- CP-element group 202: 	 assign_stmt_89_to_assign_stmt_1130/slice_278_Sample/ra
      -- 
    ra_1235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_278_inst_ack_0, ack => maxPool4_CP_307_elements(202)); -- 
    -- CP-element group 203:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	201 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	338 
    -- CP-element group 203: marked-successors 
    -- CP-element group 203: 	201 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 assign_stmt_89_to_assign_stmt_1130/slice_278_update_completed_
      -- CP-element group 203: 	 assign_stmt_89_to_assign_stmt_1130/slice_278_Update/$exit
      -- CP-element group 203: 	 assign_stmt_89_to_assign_stmt_1130/slice_278_Update/ca
      -- 
    ca_1240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_278_inst_ack_1, ack => maxPool4_CP_307_elements(203)); -- 
    -- CP-element group 204:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	47 
    -- CP-element group 204: marked-predecessors 
    -- CP-element group 204: 	206 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	206 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 assign_stmt_89_to_assign_stmt_1130/slice_282_sample_start_
      -- CP-element group 204: 	 assign_stmt_89_to_assign_stmt_1130/slice_282_Sample/$entry
      -- CP-element group 204: 	 assign_stmt_89_to_assign_stmt_1130/slice_282_Sample/rr
      -- 
    rr_1248_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1248_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(204), ack => slice_282_inst_req_0); -- 
    maxPool4_cp_element_group_204: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_204"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(47) & maxPool4_CP_307_elements(206);
      gj_maxPool4_cp_element_group_204 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(204), clk => clk, reset => reset); --
    end block;
    -- CP-element group 205:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: marked-predecessors 
    -- CP-element group 205: 	207 
    -- CP-element group 205: 	340 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	207 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 assign_stmt_89_to_assign_stmt_1130/slice_282_update_start_
      -- CP-element group 205: 	 assign_stmt_89_to_assign_stmt_1130/slice_282_Update/$entry
      -- CP-element group 205: 	 assign_stmt_89_to_assign_stmt_1130/slice_282_Update/cr
      -- 
    cr_1253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(205), ack => slice_282_inst_req_1); -- 
    maxPool4_cp_element_group_205: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_205"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(207) & maxPool4_CP_307_elements(340);
      gj_maxPool4_cp_element_group_205 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(205), clk => clk, reset => reset); --
    end block;
    -- CP-element group 206:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	204 
    -- CP-element group 206: successors 
    -- CP-element group 206: marked-successors 
    -- CP-element group 206: 	45 
    -- CP-element group 206: 	204 
    -- CP-element group 206:  members (3) 
      -- CP-element group 206: 	 assign_stmt_89_to_assign_stmt_1130/slice_282_sample_completed_
      -- CP-element group 206: 	 assign_stmt_89_to_assign_stmt_1130/slice_282_Sample/$exit
      -- CP-element group 206: 	 assign_stmt_89_to_assign_stmt_1130/slice_282_Sample/ra
      -- 
    ra_1249_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_282_inst_ack_0, ack => maxPool4_CP_307_elements(206)); -- 
    -- CP-element group 207:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	205 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	338 
    -- CP-element group 207: marked-successors 
    -- CP-element group 207: 	205 
    -- CP-element group 207:  members (3) 
      -- CP-element group 207: 	 assign_stmt_89_to_assign_stmt_1130/slice_282_update_completed_
      -- CP-element group 207: 	 assign_stmt_89_to_assign_stmt_1130/slice_282_Update/$exit
      -- CP-element group 207: 	 assign_stmt_89_to_assign_stmt_1130/slice_282_Update/ca
      -- 
    ca_1254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_282_inst_ack_1, ack => maxPool4_CP_307_elements(207)); -- 
    -- CP-element group 208:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	47 
    -- CP-element group 208: marked-predecessors 
    -- CP-element group 208: 	210 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	210 
    -- CP-element group 208:  members (3) 
      -- CP-element group 208: 	 assign_stmt_89_to_assign_stmt_1130/slice_286_sample_start_
      -- CP-element group 208: 	 assign_stmt_89_to_assign_stmt_1130/slice_286_Sample/$entry
      -- CP-element group 208: 	 assign_stmt_89_to_assign_stmt_1130/slice_286_Sample/rr
      -- 
    rr_1262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(208), ack => slice_286_inst_req_0); -- 
    maxPool4_cp_element_group_208: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_208"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(47) & maxPool4_CP_307_elements(210);
      gj_maxPool4_cp_element_group_208 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(208), clk => clk, reset => reset); --
    end block;
    -- CP-element group 209:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: marked-predecessors 
    -- CP-element group 209: 	211 
    -- CP-element group 209: 	340 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	211 
    -- CP-element group 209:  members (3) 
      -- CP-element group 209: 	 assign_stmt_89_to_assign_stmt_1130/slice_286_update_start_
      -- CP-element group 209: 	 assign_stmt_89_to_assign_stmt_1130/slice_286_Update/$entry
      -- CP-element group 209: 	 assign_stmt_89_to_assign_stmt_1130/slice_286_Update/cr
      -- 
    cr_1267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(209), ack => slice_286_inst_req_1); -- 
    maxPool4_cp_element_group_209: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_209"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(211) & maxPool4_CP_307_elements(340);
      gj_maxPool4_cp_element_group_209 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(209), clk => clk, reset => reset); --
    end block;
    -- CP-element group 210:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	208 
    -- CP-element group 210: successors 
    -- CP-element group 210: marked-successors 
    -- CP-element group 210: 	45 
    -- CP-element group 210: 	208 
    -- CP-element group 210:  members (3) 
      -- CP-element group 210: 	 assign_stmt_89_to_assign_stmt_1130/slice_286_sample_completed_
      -- CP-element group 210: 	 assign_stmt_89_to_assign_stmt_1130/slice_286_Sample/$exit
      -- CP-element group 210: 	 assign_stmt_89_to_assign_stmt_1130/slice_286_Sample/ra
      -- 
    ra_1263_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_286_inst_ack_0, ack => maxPool4_CP_307_elements(210)); -- 
    -- CP-element group 211:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	209 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	338 
    -- CP-element group 211: marked-successors 
    -- CP-element group 211: 	209 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 assign_stmt_89_to_assign_stmt_1130/slice_286_update_completed_
      -- CP-element group 211: 	 assign_stmt_89_to_assign_stmt_1130/slice_286_Update/$exit
      -- CP-element group 211: 	 assign_stmt_89_to_assign_stmt_1130/slice_286_Update/ca
      -- 
    ca_1268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_286_inst_ack_1, ack => maxPool4_CP_307_elements(211)); -- 
    -- CP-element group 212:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	47 
    -- CP-element group 212: marked-predecessors 
    -- CP-element group 212: 	214 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	214 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 assign_stmt_89_to_assign_stmt_1130/slice_290_sample_start_
      -- CP-element group 212: 	 assign_stmt_89_to_assign_stmt_1130/slice_290_Sample/$entry
      -- CP-element group 212: 	 assign_stmt_89_to_assign_stmt_1130/slice_290_Sample/rr
      -- 
    rr_1276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(212), ack => slice_290_inst_req_0); -- 
    maxPool4_cp_element_group_212: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_212"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(47) & maxPool4_CP_307_elements(214);
      gj_maxPool4_cp_element_group_212 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(212), clk => clk, reset => reset); --
    end block;
    -- CP-element group 213:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: marked-predecessors 
    -- CP-element group 213: 	215 
    -- CP-element group 213: 	359 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	215 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 assign_stmt_89_to_assign_stmt_1130/slice_290_update_start_
      -- CP-element group 213: 	 assign_stmt_89_to_assign_stmt_1130/slice_290_Update/$entry
      -- CP-element group 213: 	 assign_stmt_89_to_assign_stmt_1130/slice_290_Update/cr
      -- 
    cr_1281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(213), ack => slice_290_inst_req_1); -- 
    maxPool4_cp_element_group_213: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_213"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(215) & maxPool4_CP_307_elements(359);
      gj_maxPool4_cp_element_group_213 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(213), clk => clk, reset => reset); --
    end block;
    -- CP-element group 214:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	212 
    -- CP-element group 214: successors 
    -- CP-element group 214: marked-successors 
    -- CP-element group 214: 	45 
    -- CP-element group 214: 	212 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 assign_stmt_89_to_assign_stmt_1130/slice_290_sample_completed_
      -- CP-element group 214: 	 assign_stmt_89_to_assign_stmt_1130/slice_290_Sample/$exit
      -- CP-element group 214: 	 assign_stmt_89_to_assign_stmt_1130/slice_290_Sample/ra
      -- 
    ra_1277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_290_inst_ack_0, ack => maxPool4_CP_307_elements(214)); -- 
    -- CP-element group 215:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	213 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	357 
    -- CP-element group 215: marked-successors 
    -- CP-element group 215: 	213 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 assign_stmt_89_to_assign_stmt_1130/slice_290_update_completed_
      -- CP-element group 215: 	 assign_stmt_89_to_assign_stmt_1130/slice_290_Update/$exit
      -- CP-element group 215: 	 assign_stmt_89_to_assign_stmt_1130/slice_290_Update/ca
      -- 
    ca_1282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_290_inst_ack_1, ack => maxPool4_CP_307_elements(215)); -- 
    -- CP-element group 216:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	47 
    -- CP-element group 216: marked-predecessors 
    -- CP-element group 216: 	218 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	218 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 assign_stmt_89_to_assign_stmt_1130/slice_294_sample_start_
      -- CP-element group 216: 	 assign_stmt_89_to_assign_stmt_1130/slice_294_Sample/$entry
      -- CP-element group 216: 	 assign_stmt_89_to_assign_stmt_1130/slice_294_Sample/rr
      -- 
    rr_1290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(216), ack => slice_294_inst_req_0); -- 
    maxPool4_cp_element_group_216: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_216"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(47) & maxPool4_CP_307_elements(218);
      gj_maxPool4_cp_element_group_216 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(216), clk => clk, reset => reset); --
    end block;
    -- CP-element group 217:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: marked-predecessors 
    -- CP-element group 217: 	219 
    -- CP-element group 217: 	359 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	219 
    -- CP-element group 217:  members (3) 
      -- CP-element group 217: 	 assign_stmt_89_to_assign_stmt_1130/slice_294_update_start_
      -- CP-element group 217: 	 assign_stmt_89_to_assign_stmt_1130/slice_294_Update/$entry
      -- CP-element group 217: 	 assign_stmt_89_to_assign_stmt_1130/slice_294_Update/cr
      -- 
    cr_1295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(217), ack => slice_294_inst_req_1); -- 
    maxPool4_cp_element_group_217: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_217"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(219) & maxPool4_CP_307_elements(359);
      gj_maxPool4_cp_element_group_217 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(217), clk => clk, reset => reset); --
    end block;
    -- CP-element group 218:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	216 
    -- CP-element group 218: successors 
    -- CP-element group 218: marked-successors 
    -- CP-element group 218: 	45 
    -- CP-element group 218: 	216 
    -- CP-element group 218:  members (3) 
      -- CP-element group 218: 	 assign_stmt_89_to_assign_stmt_1130/slice_294_sample_completed_
      -- CP-element group 218: 	 assign_stmt_89_to_assign_stmt_1130/slice_294_Sample/$exit
      -- CP-element group 218: 	 assign_stmt_89_to_assign_stmt_1130/slice_294_Sample/ra
      -- 
    ra_1291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_294_inst_ack_0, ack => maxPool4_CP_307_elements(218)); -- 
    -- CP-element group 219:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	217 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	357 
    -- CP-element group 219: marked-successors 
    -- CP-element group 219: 	217 
    -- CP-element group 219:  members (3) 
      -- CP-element group 219: 	 assign_stmt_89_to_assign_stmt_1130/slice_294_update_completed_
      -- CP-element group 219: 	 assign_stmt_89_to_assign_stmt_1130/slice_294_Update/$exit
      -- CP-element group 219: 	 assign_stmt_89_to_assign_stmt_1130/slice_294_Update/ca
      -- 
    ca_1296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_294_inst_ack_1, ack => maxPool4_CP_307_elements(219)); -- 
    -- CP-element group 220:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	47 
    -- CP-element group 220: marked-predecessors 
    -- CP-element group 220: 	222 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	222 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 assign_stmt_89_to_assign_stmt_1130/slice_298_sample_start_
      -- CP-element group 220: 	 assign_stmt_89_to_assign_stmt_1130/slice_298_Sample/$entry
      -- CP-element group 220: 	 assign_stmt_89_to_assign_stmt_1130/slice_298_Sample/rr
      -- 
    rr_1304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(220), ack => slice_298_inst_req_0); -- 
    maxPool4_cp_element_group_220: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_220"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(47) & maxPool4_CP_307_elements(222);
      gj_maxPool4_cp_element_group_220 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(220), clk => clk, reset => reset); --
    end block;
    -- CP-element group 221:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: marked-predecessors 
    -- CP-element group 221: 	223 
    -- CP-element group 221: 	359 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	223 
    -- CP-element group 221:  members (3) 
      -- CP-element group 221: 	 assign_stmt_89_to_assign_stmt_1130/slice_298_update_start_
      -- CP-element group 221: 	 assign_stmt_89_to_assign_stmt_1130/slice_298_Update/$entry
      -- CP-element group 221: 	 assign_stmt_89_to_assign_stmt_1130/slice_298_Update/cr
      -- 
    cr_1309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(221), ack => slice_298_inst_req_1); -- 
    maxPool4_cp_element_group_221: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_221"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(223) & maxPool4_CP_307_elements(359);
      gj_maxPool4_cp_element_group_221 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(221), clk => clk, reset => reset); --
    end block;
    -- CP-element group 222:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	220 
    -- CP-element group 222: successors 
    -- CP-element group 222: marked-successors 
    -- CP-element group 222: 	45 
    -- CP-element group 222: 	220 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 assign_stmt_89_to_assign_stmt_1130/slice_298_sample_completed_
      -- CP-element group 222: 	 assign_stmt_89_to_assign_stmt_1130/slice_298_Sample/$exit
      -- CP-element group 222: 	 assign_stmt_89_to_assign_stmt_1130/slice_298_Sample/ra
      -- 
    ra_1305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_298_inst_ack_0, ack => maxPool4_CP_307_elements(222)); -- 
    -- CP-element group 223:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	221 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	357 
    -- CP-element group 223: marked-successors 
    -- CP-element group 223: 	221 
    -- CP-element group 223:  members (3) 
      -- CP-element group 223: 	 assign_stmt_89_to_assign_stmt_1130/slice_298_update_completed_
      -- CP-element group 223: 	 assign_stmt_89_to_assign_stmt_1130/slice_298_Update/$exit
      -- CP-element group 223: 	 assign_stmt_89_to_assign_stmt_1130/slice_298_Update/ca
      -- 
    ca_1310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_298_inst_ack_1, ack => maxPool4_CP_307_elements(223)); -- 
    -- CP-element group 224:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	47 
    -- CP-element group 224: marked-predecessors 
    -- CP-element group 224: 	226 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	226 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 assign_stmt_89_to_assign_stmt_1130/slice_302_sample_start_
      -- CP-element group 224: 	 assign_stmt_89_to_assign_stmt_1130/slice_302_Sample/$entry
      -- CP-element group 224: 	 assign_stmt_89_to_assign_stmt_1130/slice_302_Sample/rr
      -- 
    rr_1318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(224), ack => slice_302_inst_req_0); -- 
    maxPool4_cp_element_group_224: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_224"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(47) & maxPool4_CP_307_elements(226);
      gj_maxPool4_cp_element_group_224 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(224), clk => clk, reset => reset); --
    end block;
    -- CP-element group 225:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: marked-predecessors 
    -- CP-element group 225: 	227 
    -- CP-element group 225: 	359 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	227 
    -- CP-element group 225:  members (3) 
      -- CP-element group 225: 	 assign_stmt_89_to_assign_stmt_1130/slice_302_update_start_
      -- CP-element group 225: 	 assign_stmt_89_to_assign_stmt_1130/slice_302_Update/$entry
      -- CP-element group 225: 	 assign_stmt_89_to_assign_stmt_1130/slice_302_Update/cr
      -- 
    cr_1323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(225), ack => slice_302_inst_req_1); -- 
    maxPool4_cp_element_group_225: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_225"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(227) & maxPool4_CP_307_elements(359);
      gj_maxPool4_cp_element_group_225 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(225), clk => clk, reset => reset); --
    end block;
    -- CP-element group 226:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	224 
    -- CP-element group 226: successors 
    -- CP-element group 226: marked-successors 
    -- CP-element group 226: 	45 
    -- CP-element group 226: 	224 
    -- CP-element group 226:  members (3) 
      -- CP-element group 226: 	 assign_stmt_89_to_assign_stmt_1130/slice_302_sample_completed_
      -- CP-element group 226: 	 assign_stmt_89_to_assign_stmt_1130/slice_302_Sample/$exit
      -- CP-element group 226: 	 assign_stmt_89_to_assign_stmt_1130/slice_302_Sample/ra
      -- 
    ra_1319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_302_inst_ack_0, ack => maxPool4_CP_307_elements(226)); -- 
    -- CP-element group 227:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	225 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	357 
    -- CP-element group 227: marked-successors 
    -- CP-element group 227: 	225 
    -- CP-element group 227:  members (3) 
      -- CP-element group 227: 	 assign_stmt_89_to_assign_stmt_1130/slice_302_update_completed_
      -- CP-element group 227: 	 assign_stmt_89_to_assign_stmt_1130/slice_302_Update/$exit
      -- CP-element group 227: 	 assign_stmt_89_to_assign_stmt_1130/slice_302_Update/ca
      -- 
    ca_1324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_302_inst_ack_1, ack => maxPool4_CP_307_elements(227)); -- 
    -- CP-element group 228:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	47 
    -- CP-element group 228: marked-predecessors 
    -- CP-element group 228: 	230 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	230 
    -- CP-element group 228:  members (3) 
      -- CP-element group 228: 	 assign_stmt_89_to_assign_stmt_1130/slice_306_sample_start_
      -- CP-element group 228: 	 assign_stmt_89_to_assign_stmt_1130/slice_306_Sample/$entry
      -- CP-element group 228: 	 assign_stmt_89_to_assign_stmt_1130/slice_306_Sample/rr
      -- 
    rr_1332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(228), ack => slice_306_inst_req_0); -- 
    maxPool4_cp_element_group_228: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_228"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(47) & maxPool4_CP_307_elements(230);
      gj_maxPool4_cp_element_group_228 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(228), clk => clk, reset => reset); --
    end block;
    -- CP-element group 229:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: marked-predecessors 
    -- CP-element group 229: 	231 
    -- CP-element group 229: 	378 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	231 
    -- CP-element group 229:  members (3) 
      -- CP-element group 229: 	 assign_stmt_89_to_assign_stmt_1130/slice_306_update_start_
      -- CP-element group 229: 	 assign_stmt_89_to_assign_stmt_1130/slice_306_Update/$entry
      -- CP-element group 229: 	 assign_stmt_89_to_assign_stmt_1130/slice_306_Update/cr
      -- 
    cr_1337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(229), ack => slice_306_inst_req_1); -- 
    maxPool4_cp_element_group_229: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_229"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(231) & maxPool4_CP_307_elements(378);
      gj_maxPool4_cp_element_group_229 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(229), clk => clk, reset => reset); --
    end block;
    -- CP-element group 230:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	228 
    -- CP-element group 230: successors 
    -- CP-element group 230: marked-successors 
    -- CP-element group 230: 	45 
    -- CP-element group 230: 	228 
    -- CP-element group 230:  members (3) 
      -- CP-element group 230: 	 assign_stmt_89_to_assign_stmt_1130/slice_306_sample_completed_
      -- CP-element group 230: 	 assign_stmt_89_to_assign_stmt_1130/slice_306_Sample/$exit
      -- CP-element group 230: 	 assign_stmt_89_to_assign_stmt_1130/slice_306_Sample/ra
      -- 
    ra_1333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_306_inst_ack_0, ack => maxPool4_CP_307_elements(230)); -- 
    -- CP-element group 231:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	229 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	376 
    -- CP-element group 231: marked-successors 
    -- CP-element group 231: 	229 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 assign_stmt_89_to_assign_stmt_1130/slice_306_update_completed_
      -- CP-element group 231: 	 assign_stmt_89_to_assign_stmt_1130/slice_306_Update/$exit
      -- CP-element group 231: 	 assign_stmt_89_to_assign_stmt_1130/slice_306_Update/ca
      -- 
    ca_1338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_306_inst_ack_1, ack => maxPool4_CP_307_elements(231)); -- 
    -- CP-element group 232:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	47 
    -- CP-element group 232: marked-predecessors 
    -- CP-element group 232: 	234 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	234 
    -- CP-element group 232:  members (3) 
      -- CP-element group 232: 	 assign_stmt_89_to_assign_stmt_1130/slice_310_sample_start_
      -- CP-element group 232: 	 assign_stmt_89_to_assign_stmt_1130/slice_310_Sample/$entry
      -- CP-element group 232: 	 assign_stmt_89_to_assign_stmt_1130/slice_310_Sample/rr
      -- 
    rr_1346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(232), ack => slice_310_inst_req_0); -- 
    maxPool4_cp_element_group_232: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_232"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(47) & maxPool4_CP_307_elements(234);
      gj_maxPool4_cp_element_group_232 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(232), clk => clk, reset => reset); --
    end block;
    -- CP-element group 233:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: marked-predecessors 
    -- CP-element group 233: 	235 
    -- CP-element group 233: 	378 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	235 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 assign_stmt_89_to_assign_stmt_1130/slice_310_update_start_
      -- CP-element group 233: 	 assign_stmt_89_to_assign_stmt_1130/slice_310_Update/$entry
      -- CP-element group 233: 	 assign_stmt_89_to_assign_stmt_1130/slice_310_Update/cr
      -- 
    cr_1351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(233), ack => slice_310_inst_req_1); -- 
    maxPool4_cp_element_group_233: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_233"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(235) & maxPool4_CP_307_elements(378);
      gj_maxPool4_cp_element_group_233 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(233), clk => clk, reset => reset); --
    end block;
    -- CP-element group 234:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	232 
    -- CP-element group 234: successors 
    -- CP-element group 234: marked-successors 
    -- CP-element group 234: 	45 
    -- CP-element group 234: 	232 
    -- CP-element group 234:  members (3) 
      -- CP-element group 234: 	 assign_stmt_89_to_assign_stmt_1130/slice_310_sample_completed_
      -- CP-element group 234: 	 assign_stmt_89_to_assign_stmt_1130/slice_310_Sample/$exit
      -- CP-element group 234: 	 assign_stmt_89_to_assign_stmt_1130/slice_310_Sample/ra
      -- 
    ra_1347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_310_inst_ack_0, ack => maxPool4_CP_307_elements(234)); -- 
    -- CP-element group 235:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	233 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	376 
    -- CP-element group 235: marked-successors 
    -- CP-element group 235: 	233 
    -- CP-element group 235:  members (3) 
      -- CP-element group 235: 	 assign_stmt_89_to_assign_stmt_1130/slice_310_update_completed_
      -- CP-element group 235: 	 assign_stmt_89_to_assign_stmt_1130/slice_310_Update/$exit
      -- CP-element group 235: 	 assign_stmt_89_to_assign_stmt_1130/slice_310_Update/ca
      -- 
    ca_1352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_310_inst_ack_1, ack => maxPool4_CP_307_elements(235)); -- 
    -- CP-element group 236:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	47 
    -- CP-element group 236: marked-predecessors 
    -- CP-element group 236: 	238 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	238 
    -- CP-element group 236:  members (3) 
      -- CP-element group 236: 	 assign_stmt_89_to_assign_stmt_1130/slice_314_sample_start_
      -- CP-element group 236: 	 assign_stmt_89_to_assign_stmt_1130/slice_314_Sample/$entry
      -- CP-element group 236: 	 assign_stmt_89_to_assign_stmt_1130/slice_314_Sample/rr
      -- 
    rr_1360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(236), ack => slice_314_inst_req_0); -- 
    maxPool4_cp_element_group_236: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_236"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(47) & maxPool4_CP_307_elements(238);
      gj_maxPool4_cp_element_group_236 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(236), clk => clk, reset => reset); --
    end block;
    -- CP-element group 237:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: marked-predecessors 
    -- CP-element group 237: 	239 
    -- CP-element group 237: 	378 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	239 
    -- CP-element group 237:  members (3) 
      -- CP-element group 237: 	 assign_stmt_89_to_assign_stmt_1130/slice_314_update_start_
      -- CP-element group 237: 	 assign_stmt_89_to_assign_stmt_1130/slice_314_Update/$entry
      -- CP-element group 237: 	 assign_stmt_89_to_assign_stmt_1130/slice_314_Update/cr
      -- 
    cr_1365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(237), ack => slice_314_inst_req_1); -- 
    maxPool4_cp_element_group_237: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_237"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(239) & maxPool4_CP_307_elements(378);
      gj_maxPool4_cp_element_group_237 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(237), clk => clk, reset => reset); --
    end block;
    -- CP-element group 238:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	236 
    -- CP-element group 238: successors 
    -- CP-element group 238: marked-successors 
    -- CP-element group 238: 	45 
    -- CP-element group 238: 	236 
    -- CP-element group 238:  members (3) 
      -- CP-element group 238: 	 assign_stmt_89_to_assign_stmt_1130/slice_314_sample_completed_
      -- CP-element group 238: 	 assign_stmt_89_to_assign_stmt_1130/slice_314_Sample/$exit
      -- CP-element group 238: 	 assign_stmt_89_to_assign_stmt_1130/slice_314_Sample/ra
      -- 
    ra_1361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_314_inst_ack_0, ack => maxPool4_CP_307_elements(238)); -- 
    -- CP-element group 239:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	237 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	376 
    -- CP-element group 239: marked-successors 
    -- CP-element group 239: 	237 
    -- CP-element group 239:  members (3) 
      -- CP-element group 239: 	 assign_stmt_89_to_assign_stmt_1130/slice_314_update_completed_
      -- CP-element group 239: 	 assign_stmt_89_to_assign_stmt_1130/slice_314_Update/$exit
      -- CP-element group 239: 	 assign_stmt_89_to_assign_stmt_1130/slice_314_Update/ca
      -- 
    ca_1366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_314_inst_ack_1, ack => maxPool4_CP_307_elements(239)); -- 
    -- CP-element group 240:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	47 
    -- CP-element group 240: marked-predecessors 
    -- CP-element group 240: 	242 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	242 
    -- CP-element group 240:  members (3) 
      -- CP-element group 240: 	 assign_stmt_89_to_assign_stmt_1130/slice_318_sample_start_
      -- CP-element group 240: 	 assign_stmt_89_to_assign_stmt_1130/slice_318_Sample/$entry
      -- CP-element group 240: 	 assign_stmt_89_to_assign_stmt_1130/slice_318_Sample/rr
      -- 
    rr_1374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(240), ack => slice_318_inst_req_0); -- 
    maxPool4_cp_element_group_240: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_240"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(47) & maxPool4_CP_307_elements(242);
      gj_maxPool4_cp_element_group_240 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(240), clk => clk, reset => reset); --
    end block;
    -- CP-element group 241:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: marked-predecessors 
    -- CP-element group 241: 	243 
    -- CP-element group 241: 	378 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	243 
    -- CP-element group 241:  members (3) 
      -- CP-element group 241: 	 assign_stmt_89_to_assign_stmt_1130/slice_318_update_start_
      -- CP-element group 241: 	 assign_stmt_89_to_assign_stmt_1130/slice_318_Update/$entry
      -- CP-element group 241: 	 assign_stmt_89_to_assign_stmt_1130/slice_318_Update/cr
      -- 
    cr_1379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(241), ack => slice_318_inst_req_1); -- 
    maxPool4_cp_element_group_241: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_241"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(243) & maxPool4_CP_307_elements(378);
      gj_maxPool4_cp_element_group_241 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(241), clk => clk, reset => reset); --
    end block;
    -- CP-element group 242:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	240 
    -- CP-element group 242: successors 
    -- CP-element group 242: marked-successors 
    -- CP-element group 242: 	45 
    -- CP-element group 242: 	240 
    -- CP-element group 242:  members (3) 
      -- CP-element group 242: 	 assign_stmt_89_to_assign_stmt_1130/slice_318_sample_completed_
      -- CP-element group 242: 	 assign_stmt_89_to_assign_stmt_1130/slice_318_Sample/$exit
      -- CP-element group 242: 	 assign_stmt_89_to_assign_stmt_1130/slice_318_Sample/ra
      -- 
    ra_1375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_318_inst_ack_0, ack => maxPool4_CP_307_elements(242)); -- 
    -- CP-element group 243:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	241 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	376 
    -- CP-element group 243: marked-successors 
    -- CP-element group 243: 	241 
    -- CP-element group 243:  members (3) 
      -- CP-element group 243: 	 assign_stmt_89_to_assign_stmt_1130/slice_318_update_completed_
      -- CP-element group 243: 	 assign_stmt_89_to_assign_stmt_1130/slice_318_Update/$exit
      -- CP-element group 243: 	 assign_stmt_89_to_assign_stmt_1130/slice_318_Update/ca
      -- 
    ca_1380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_318_inst_ack_1, ack => maxPool4_CP_307_elements(243)); -- 
    -- CP-element group 244:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	51 
    -- CP-element group 244: marked-predecessors 
    -- CP-element group 244: 	246 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	246 
    -- CP-element group 244:  members (3) 
      -- CP-element group 244: 	 assign_stmt_89_to_assign_stmt_1130/slice_322_sample_start_
      -- CP-element group 244: 	 assign_stmt_89_to_assign_stmt_1130/slice_322_Sample/$entry
      -- CP-element group 244: 	 assign_stmt_89_to_assign_stmt_1130/slice_322_Sample/rr
      -- 
    rr_1388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(244), ack => slice_322_inst_req_0); -- 
    maxPool4_cp_element_group_244: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_244"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(51) & maxPool4_CP_307_elements(246);
      gj_maxPool4_cp_element_group_244 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(244), clk => clk, reset => reset); --
    end block;
    -- CP-element group 245:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: marked-predecessors 
    -- CP-element group 245: 	247 
    -- CP-element group 245: 	321 
    -- CP-element group 245: 	386 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	247 
    -- CP-element group 245:  members (3) 
      -- CP-element group 245: 	 assign_stmt_89_to_assign_stmt_1130/slice_322_update_start_
      -- CP-element group 245: 	 assign_stmt_89_to_assign_stmt_1130/slice_322_Update/$entry
      -- CP-element group 245: 	 assign_stmt_89_to_assign_stmt_1130/slice_322_Update/cr
      -- 
    cr_1393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(245), ack => slice_322_inst_req_1); -- 
    maxPool4_cp_element_group_245: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_245"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(247) & maxPool4_CP_307_elements(321) & maxPool4_CP_307_elements(386);
      gj_maxPool4_cp_element_group_245 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(245), clk => clk, reset => reset); --
    end block;
    -- CP-element group 246:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	244 
    -- CP-element group 246: successors 
    -- CP-element group 246: marked-successors 
    -- CP-element group 246: 	49 
    -- CP-element group 246: 	244 
    -- CP-element group 246:  members (3) 
      -- CP-element group 246: 	 assign_stmt_89_to_assign_stmt_1130/slice_322_sample_completed_
      -- CP-element group 246: 	 assign_stmt_89_to_assign_stmt_1130/slice_322_Sample/$exit
      -- CP-element group 246: 	 assign_stmt_89_to_assign_stmt_1130/slice_322_Sample/ra
      -- 
    ra_1389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_322_inst_ack_0, ack => maxPool4_CP_307_elements(246)); -- 
    -- CP-element group 247:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	245 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	319 
    -- CP-element group 247: 	384 
    -- CP-element group 247: marked-successors 
    -- CP-element group 247: 	245 
    -- CP-element group 247:  members (3) 
      -- CP-element group 247: 	 assign_stmt_89_to_assign_stmt_1130/slice_322_update_completed_
      -- CP-element group 247: 	 assign_stmt_89_to_assign_stmt_1130/slice_322_Update/$exit
      -- CP-element group 247: 	 assign_stmt_89_to_assign_stmt_1130/slice_322_Update/ca
      -- 
    ca_1394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_322_inst_ack_1, ack => maxPool4_CP_307_elements(247)); -- 
    -- CP-element group 248:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	51 
    -- CP-element group 248: marked-predecessors 
    -- CP-element group 248: 	250 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	250 
    -- CP-element group 248:  members (3) 
      -- CP-element group 248: 	 assign_stmt_89_to_assign_stmt_1130/slice_326_sample_start_
      -- CP-element group 248: 	 assign_stmt_89_to_assign_stmt_1130/slice_326_Sample/$entry
      -- CP-element group 248: 	 assign_stmt_89_to_assign_stmt_1130/slice_326_Sample/rr
      -- 
    rr_1402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(248), ack => slice_326_inst_req_0); -- 
    maxPool4_cp_element_group_248: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_248"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(51) & maxPool4_CP_307_elements(250);
      gj_maxPool4_cp_element_group_248 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(248), clk => clk, reset => reset); --
    end block;
    -- CP-element group 249:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: marked-predecessors 
    -- CP-element group 249: 	251 
    -- CP-element group 249: 	321 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	251 
    -- CP-element group 249:  members (3) 
      -- CP-element group 249: 	 assign_stmt_89_to_assign_stmt_1130/slice_326_update_start_
      -- CP-element group 249: 	 assign_stmt_89_to_assign_stmt_1130/slice_326_Update/$entry
      -- CP-element group 249: 	 assign_stmt_89_to_assign_stmt_1130/slice_326_Update/cr
      -- 
    cr_1407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(249), ack => slice_326_inst_req_1); -- 
    maxPool4_cp_element_group_249: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_249"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(251) & maxPool4_CP_307_elements(321);
      gj_maxPool4_cp_element_group_249 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(249), clk => clk, reset => reset); --
    end block;
    -- CP-element group 250:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	248 
    -- CP-element group 250: successors 
    -- CP-element group 250: marked-successors 
    -- CP-element group 250: 	49 
    -- CP-element group 250: 	248 
    -- CP-element group 250:  members (3) 
      -- CP-element group 250: 	 assign_stmt_89_to_assign_stmt_1130/slice_326_sample_completed_
      -- CP-element group 250: 	 assign_stmt_89_to_assign_stmt_1130/slice_326_Sample/$exit
      -- CP-element group 250: 	 assign_stmt_89_to_assign_stmt_1130/slice_326_Sample/ra
      -- 
    ra_1403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_326_inst_ack_0, ack => maxPool4_CP_307_elements(250)); -- 
    -- CP-element group 251:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	249 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	319 
    -- CP-element group 251: marked-successors 
    -- CP-element group 251: 	249 
    -- CP-element group 251:  members (3) 
      -- CP-element group 251: 	 assign_stmt_89_to_assign_stmt_1130/slice_326_update_completed_
      -- CP-element group 251: 	 assign_stmt_89_to_assign_stmt_1130/slice_326_Update/$exit
      -- CP-element group 251: 	 assign_stmt_89_to_assign_stmt_1130/slice_326_Update/ca
      -- 
    ca_1408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_326_inst_ack_1, ack => maxPool4_CP_307_elements(251)); -- 
    -- CP-element group 252:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	51 
    -- CP-element group 252: marked-predecessors 
    -- CP-element group 252: 	254 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	254 
    -- CP-element group 252:  members (3) 
      -- CP-element group 252: 	 assign_stmt_89_to_assign_stmt_1130/slice_330_sample_start_
      -- CP-element group 252: 	 assign_stmt_89_to_assign_stmt_1130/slice_330_Sample/$entry
      -- CP-element group 252: 	 assign_stmt_89_to_assign_stmt_1130/slice_330_Sample/rr
      -- 
    rr_1416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(252), ack => slice_330_inst_req_0); -- 
    maxPool4_cp_element_group_252: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_252"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(51) & maxPool4_CP_307_elements(254);
      gj_maxPool4_cp_element_group_252 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(252), clk => clk, reset => reset); --
    end block;
    -- CP-element group 253:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: marked-predecessors 
    -- CP-element group 253: 	255 
    -- CP-element group 253: 	321 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	255 
    -- CP-element group 253:  members (3) 
      -- CP-element group 253: 	 assign_stmt_89_to_assign_stmt_1130/slice_330_update_start_
      -- CP-element group 253: 	 assign_stmt_89_to_assign_stmt_1130/slice_330_Update/$entry
      -- CP-element group 253: 	 assign_stmt_89_to_assign_stmt_1130/slice_330_Update/cr
      -- 
    cr_1421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(253), ack => slice_330_inst_req_1); -- 
    maxPool4_cp_element_group_253: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_253"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(255) & maxPool4_CP_307_elements(321);
      gj_maxPool4_cp_element_group_253 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(253), clk => clk, reset => reset); --
    end block;
    -- CP-element group 254:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	252 
    -- CP-element group 254: successors 
    -- CP-element group 254: marked-successors 
    -- CP-element group 254: 	49 
    -- CP-element group 254: 	252 
    -- CP-element group 254:  members (3) 
      -- CP-element group 254: 	 assign_stmt_89_to_assign_stmt_1130/slice_330_sample_completed_
      -- CP-element group 254: 	 assign_stmt_89_to_assign_stmt_1130/slice_330_Sample/$exit
      -- CP-element group 254: 	 assign_stmt_89_to_assign_stmt_1130/slice_330_Sample/ra
      -- 
    ra_1417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_330_inst_ack_0, ack => maxPool4_CP_307_elements(254)); -- 
    -- CP-element group 255:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	253 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	319 
    -- CP-element group 255: marked-successors 
    -- CP-element group 255: 	253 
    -- CP-element group 255:  members (3) 
      -- CP-element group 255: 	 assign_stmt_89_to_assign_stmt_1130/slice_330_update_completed_
      -- CP-element group 255: 	 assign_stmt_89_to_assign_stmt_1130/slice_330_Update/$exit
      -- CP-element group 255: 	 assign_stmt_89_to_assign_stmt_1130/slice_330_Update/ca
      -- 
    ca_1422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_330_inst_ack_1, ack => maxPool4_CP_307_elements(255)); -- 
    -- CP-element group 256:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	51 
    -- CP-element group 256: marked-predecessors 
    -- CP-element group 256: 	258 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	258 
    -- CP-element group 256:  members (3) 
      -- CP-element group 256: 	 assign_stmt_89_to_assign_stmt_1130/slice_334_sample_start_
      -- CP-element group 256: 	 assign_stmt_89_to_assign_stmt_1130/slice_334_Sample/$entry
      -- CP-element group 256: 	 assign_stmt_89_to_assign_stmt_1130/slice_334_Sample/rr
      -- 
    rr_1430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(256), ack => slice_334_inst_req_0); -- 
    maxPool4_cp_element_group_256: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_256"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(51) & maxPool4_CP_307_elements(258);
      gj_maxPool4_cp_element_group_256 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(256), clk => clk, reset => reset); --
    end block;
    -- CP-element group 257:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: marked-predecessors 
    -- CP-element group 257: 	259 
    -- CP-element group 257: 	321 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	259 
    -- CP-element group 257:  members (3) 
      -- CP-element group 257: 	 assign_stmt_89_to_assign_stmt_1130/slice_334_update_start_
      -- CP-element group 257: 	 assign_stmt_89_to_assign_stmt_1130/slice_334_Update/$entry
      -- CP-element group 257: 	 assign_stmt_89_to_assign_stmt_1130/slice_334_Update/cr
      -- 
    cr_1435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(257), ack => slice_334_inst_req_1); -- 
    maxPool4_cp_element_group_257: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_257"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(259) & maxPool4_CP_307_elements(321);
      gj_maxPool4_cp_element_group_257 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(257), clk => clk, reset => reset); --
    end block;
    -- CP-element group 258:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	256 
    -- CP-element group 258: successors 
    -- CP-element group 258: marked-successors 
    -- CP-element group 258: 	49 
    -- CP-element group 258: 	256 
    -- CP-element group 258:  members (3) 
      -- CP-element group 258: 	 assign_stmt_89_to_assign_stmt_1130/slice_334_sample_completed_
      -- CP-element group 258: 	 assign_stmt_89_to_assign_stmt_1130/slice_334_Sample/$exit
      -- CP-element group 258: 	 assign_stmt_89_to_assign_stmt_1130/slice_334_Sample/ra
      -- 
    ra_1431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_334_inst_ack_0, ack => maxPool4_CP_307_elements(258)); -- 
    -- CP-element group 259:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	257 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	319 
    -- CP-element group 259: marked-successors 
    -- CP-element group 259: 	257 
    -- CP-element group 259:  members (3) 
      -- CP-element group 259: 	 assign_stmt_89_to_assign_stmt_1130/slice_334_update_completed_
      -- CP-element group 259: 	 assign_stmt_89_to_assign_stmt_1130/slice_334_Update/$exit
      -- CP-element group 259: 	 assign_stmt_89_to_assign_stmt_1130/slice_334_Update/ca
      -- 
    ca_1436_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_334_inst_ack_1, ack => maxPool4_CP_307_elements(259)); -- 
    -- CP-element group 260:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	51 
    -- CP-element group 260: marked-predecessors 
    -- CP-element group 260: 	262 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	262 
    -- CP-element group 260:  members (3) 
      -- CP-element group 260: 	 assign_stmt_89_to_assign_stmt_1130/slice_338_sample_start_
      -- CP-element group 260: 	 assign_stmt_89_to_assign_stmt_1130/slice_338_Sample/$entry
      -- CP-element group 260: 	 assign_stmt_89_to_assign_stmt_1130/slice_338_Sample/rr
      -- 
    rr_1444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(260), ack => slice_338_inst_req_0); -- 
    maxPool4_cp_element_group_260: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_260"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(51) & maxPool4_CP_307_elements(262);
      gj_maxPool4_cp_element_group_260 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(260), clk => clk, reset => reset); --
    end block;
    -- CP-element group 261:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: marked-predecessors 
    -- CP-element group 261: 	263 
    -- CP-element group 261: 	340 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	263 
    -- CP-element group 261:  members (3) 
      -- CP-element group 261: 	 assign_stmt_89_to_assign_stmt_1130/slice_338_update_start_
      -- CP-element group 261: 	 assign_stmt_89_to_assign_stmt_1130/slice_338_Update/$entry
      -- CP-element group 261: 	 assign_stmt_89_to_assign_stmt_1130/slice_338_Update/cr
      -- 
    cr_1449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(261), ack => slice_338_inst_req_1); -- 
    maxPool4_cp_element_group_261: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_261"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(263) & maxPool4_CP_307_elements(340);
      gj_maxPool4_cp_element_group_261 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(261), clk => clk, reset => reset); --
    end block;
    -- CP-element group 262:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	260 
    -- CP-element group 262: successors 
    -- CP-element group 262: marked-successors 
    -- CP-element group 262: 	49 
    -- CP-element group 262: 	260 
    -- CP-element group 262:  members (3) 
      -- CP-element group 262: 	 assign_stmt_89_to_assign_stmt_1130/slice_338_sample_completed_
      -- CP-element group 262: 	 assign_stmt_89_to_assign_stmt_1130/slice_338_Sample/$exit
      -- CP-element group 262: 	 assign_stmt_89_to_assign_stmt_1130/slice_338_Sample/ra
      -- 
    ra_1445_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_338_inst_ack_0, ack => maxPool4_CP_307_elements(262)); -- 
    -- CP-element group 263:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	261 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	338 
    -- CP-element group 263: marked-successors 
    -- CP-element group 263: 	261 
    -- CP-element group 263:  members (3) 
      -- CP-element group 263: 	 assign_stmt_89_to_assign_stmt_1130/slice_338_update_completed_
      -- CP-element group 263: 	 assign_stmt_89_to_assign_stmt_1130/slice_338_Update/$exit
      -- CP-element group 263: 	 assign_stmt_89_to_assign_stmt_1130/slice_338_Update/ca
      -- 
    ca_1450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_338_inst_ack_1, ack => maxPool4_CP_307_elements(263)); -- 
    -- CP-element group 264:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	51 
    -- CP-element group 264: marked-predecessors 
    -- CP-element group 264: 	266 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	266 
    -- CP-element group 264:  members (3) 
      -- CP-element group 264: 	 assign_stmt_89_to_assign_stmt_1130/slice_342_sample_start_
      -- CP-element group 264: 	 assign_stmt_89_to_assign_stmt_1130/slice_342_Sample/$entry
      -- CP-element group 264: 	 assign_stmt_89_to_assign_stmt_1130/slice_342_Sample/rr
      -- 
    rr_1458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(264), ack => slice_342_inst_req_0); -- 
    maxPool4_cp_element_group_264: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_264"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(51) & maxPool4_CP_307_elements(266);
      gj_maxPool4_cp_element_group_264 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(264), clk => clk, reset => reset); --
    end block;
    -- CP-element group 265:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: marked-predecessors 
    -- CP-element group 265: 	267 
    -- CP-element group 265: 	340 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	267 
    -- CP-element group 265:  members (3) 
      -- CP-element group 265: 	 assign_stmt_89_to_assign_stmt_1130/slice_342_update_start_
      -- CP-element group 265: 	 assign_stmt_89_to_assign_stmt_1130/slice_342_Update/$entry
      -- CP-element group 265: 	 assign_stmt_89_to_assign_stmt_1130/slice_342_Update/cr
      -- 
    cr_1463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(265), ack => slice_342_inst_req_1); -- 
    maxPool4_cp_element_group_265: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_265"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(267) & maxPool4_CP_307_elements(340);
      gj_maxPool4_cp_element_group_265 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(265), clk => clk, reset => reset); --
    end block;
    -- CP-element group 266:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	264 
    -- CP-element group 266: successors 
    -- CP-element group 266: marked-successors 
    -- CP-element group 266: 	49 
    -- CP-element group 266: 	264 
    -- CP-element group 266:  members (3) 
      -- CP-element group 266: 	 assign_stmt_89_to_assign_stmt_1130/slice_342_sample_completed_
      -- CP-element group 266: 	 assign_stmt_89_to_assign_stmt_1130/slice_342_Sample/$exit
      -- CP-element group 266: 	 assign_stmt_89_to_assign_stmt_1130/slice_342_Sample/ra
      -- 
    ra_1459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_342_inst_ack_0, ack => maxPool4_CP_307_elements(266)); -- 
    -- CP-element group 267:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	265 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	338 
    -- CP-element group 267: marked-successors 
    -- CP-element group 267: 	265 
    -- CP-element group 267:  members (3) 
      -- CP-element group 267: 	 assign_stmt_89_to_assign_stmt_1130/slice_342_update_completed_
      -- CP-element group 267: 	 assign_stmt_89_to_assign_stmt_1130/slice_342_Update/$exit
      -- CP-element group 267: 	 assign_stmt_89_to_assign_stmt_1130/slice_342_Update/ca
      -- 
    ca_1464_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_342_inst_ack_1, ack => maxPool4_CP_307_elements(267)); -- 
    -- CP-element group 268:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	51 
    -- CP-element group 268: marked-predecessors 
    -- CP-element group 268: 	270 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	270 
    -- CP-element group 268:  members (3) 
      -- CP-element group 268: 	 assign_stmt_89_to_assign_stmt_1130/slice_346_sample_start_
      -- CP-element group 268: 	 assign_stmt_89_to_assign_stmt_1130/slice_346_Sample/$entry
      -- CP-element group 268: 	 assign_stmt_89_to_assign_stmt_1130/slice_346_Sample/rr
      -- 
    rr_1472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(268), ack => slice_346_inst_req_0); -- 
    maxPool4_cp_element_group_268: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_268"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(51) & maxPool4_CP_307_elements(270);
      gj_maxPool4_cp_element_group_268 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(268), clk => clk, reset => reset); --
    end block;
    -- CP-element group 269:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: marked-predecessors 
    -- CP-element group 269: 	271 
    -- CP-element group 269: 	340 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	271 
    -- CP-element group 269:  members (3) 
      -- CP-element group 269: 	 assign_stmt_89_to_assign_stmt_1130/slice_346_update_start_
      -- CP-element group 269: 	 assign_stmt_89_to_assign_stmt_1130/slice_346_Update/$entry
      -- CP-element group 269: 	 assign_stmt_89_to_assign_stmt_1130/slice_346_Update/cr
      -- 
    cr_1477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(269), ack => slice_346_inst_req_1); -- 
    maxPool4_cp_element_group_269: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_269"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(271) & maxPool4_CP_307_elements(340);
      gj_maxPool4_cp_element_group_269 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(269), clk => clk, reset => reset); --
    end block;
    -- CP-element group 270:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	268 
    -- CP-element group 270: successors 
    -- CP-element group 270: marked-successors 
    -- CP-element group 270: 	49 
    -- CP-element group 270: 	268 
    -- CP-element group 270:  members (3) 
      -- CP-element group 270: 	 assign_stmt_89_to_assign_stmt_1130/slice_346_sample_completed_
      -- CP-element group 270: 	 assign_stmt_89_to_assign_stmt_1130/slice_346_Sample/$exit
      -- CP-element group 270: 	 assign_stmt_89_to_assign_stmt_1130/slice_346_Sample/ra
      -- 
    ra_1473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_346_inst_ack_0, ack => maxPool4_CP_307_elements(270)); -- 
    -- CP-element group 271:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	269 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	338 
    -- CP-element group 271: marked-successors 
    -- CP-element group 271: 	269 
    -- CP-element group 271:  members (3) 
      -- CP-element group 271: 	 assign_stmt_89_to_assign_stmt_1130/slice_346_update_completed_
      -- CP-element group 271: 	 assign_stmt_89_to_assign_stmt_1130/slice_346_Update/$exit
      -- CP-element group 271: 	 assign_stmt_89_to_assign_stmt_1130/slice_346_Update/ca
      -- 
    ca_1478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_346_inst_ack_1, ack => maxPool4_CP_307_elements(271)); -- 
    -- CP-element group 272:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	51 
    -- CP-element group 272: marked-predecessors 
    -- CP-element group 272: 	274 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	274 
    -- CP-element group 272:  members (3) 
      -- CP-element group 272: 	 assign_stmt_89_to_assign_stmt_1130/slice_350_sample_start_
      -- CP-element group 272: 	 assign_stmt_89_to_assign_stmt_1130/slice_350_Sample/$entry
      -- CP-element group 272: 	 assign_stmt_89_to_assign_stmt_1130/slice_350_Sample/rr
      -- 
    rr_1486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(272), ack => slice_350_inst_req_0); -- 
    maxPool4_cp_element_group_272: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_272"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(51) & maxPool4_CP_307_elements(274);
      gj_maxPool4_cp_element_group_272 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(272), clk => clk, reset => reset); --
    end block;
    -- CP-element group 273:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: marked-predecessors 
    -- CP-element group 273: 	275 
    -- CP-element group 273: 	340 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	275 
    -- CP-element group 273:  members (3) 
      -- CP-element group 273: 	 assign_stmt_89_to_assign_stmt_1130/slice_350_update_start_
      -- CP-element group 273: 	 assign_stmt_89_to_assign_stmt_1130/slice_350_Update/$entry
      -- CP-element group 273: 	 assign_stmt_89_to_assign_stmt_1130/slice_350_Update/cr
      -- 
    cr_1491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(273), ack => slice_350_inst_req_1); -- 
    maxPool4_cp_element_group_273: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_273"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(275) & maxPool4_CP_307_elements(340);
      gj_maxPool4_cp_element_group_273 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(273), clk => clk, reset => reset); --
    end block;
    -- CP-element group 274:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	272 
    -- CP-element group 274: successors 
    -- CP-element group 274: marked-successors 
    -- CP-element group 274: 	49 
    -- CP-element group 274: 	272 
    -- CP-element group 274:  members (3) 
      -- CP-element group 274: 	 assign_stmt_89_to_assign_stmt_1130/slice_350_sample_completed_
      -- CP-element group 274: 	 assign_stmt_89_to_assign_stmt_1130/slice_350_Sample/$exit
      -- CP-element group 274: 	 assign_stmt_89_to_assign_stmt_1130/slice_350_Sample/ra
      -- 
    ra_1487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_350_inst_ack_0, ack => maxPool4_CP_307_elements(274)); -- 
    -- CP-element group 275:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	273 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	338 
    -- CP-element group 275: marked-successors 
    -- CP-element group 275: 	273 
    -- CP-element group 275:  members (3) 
      -- CP-element group 275: 	 assign_stmt_89_to_assign_stmt_1130/slice_350_update_completed_
      -- CP-element group 275: 	 assign_stmt_89_to_assign_stmt_1130/slice_350_Update/$exit
      -- CP-element group 275: 	 assign_stmt_89_to_assign_stmt_1130/slice_350_Update/ca
      -- 
    ca_1492_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_350_inst_ack_1, ack => maxPool4_CP_307_elements(275)); -- 
    -- CP-element group 276:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	51 
    -- CP-element group 276: marked-predecessors 
    -- CP-element group 276: 	278 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	278 
    -- CP-element group 276:  members (3) 
      -- CP-element group 276: 	 assign_stmt_89_to_assign_stmt_1130/slice_354_sample_start_
      -- CP-element group 276: 	 assign_stmt_89_to_assign_stmt_1130/slice_354_Sample/$entry
      -- CP-element group 276: 	 assign_stmt_89_to_assign_stmt_1130/slice_354_Sample/rr
      -- 
    rr_1500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(276), ack => slice_354_inst_req_0); -- 
    maxPool4_cp_element_group_276: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_276"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(51) & maxPool4_CP_307_elements(278);
      gj_maxPool4_cp_element_group_276 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(276), clk => clk, reset => reset); --
    end block;
    -- CP-element group 277:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: marked-predecessors 
    -- CP-element group 277: 	279 
    -- CP-element group 277: 	359 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	279 
    -- CP-element group 277:  members (3) 
      -- CP-element group 277: 	 assign_stmt_89_to_assign_stmt_1130/slice_354_update_start_
      -- CP-element group 277: 	 assign_stmt_89_to_assign_stmt_1130/slice_354_Update/$entry
      -- CP-element group 277: 	 assign_stmt_89_to_assign_stmt_1130/slice_354_Update/cr
      -- 
    cr_1505_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1505_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(277), ack => slice_354_inst_req_1); -- 
    maxPool4_cp_element_group_277: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_277"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(279) & maxPool4_CP_307_elements(359);
      gj_maxPool4_cp_element_group_277 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(277), clk => clk, reset => reset); --
    end block;
    -- CP-element group 278:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	276 
    -- CP-element group 278: successors 
    -- CP-element group 278: marked-successors 
    -- CP-element group 278: 	49 
    -- CP-element group 278: 	276 
    -- CP-element group 278:  members (3) 
      -- CP-element group 278: 	 assign_stmt_89_to_assign_stmt_1130/slice_354_sample_completed_
      -- CP-element group 278: 	 assign_stmt_89_to_assign_stmt_1130/slice_354_Sample/$exit
      -- CP-element group 278: 	 assign_stmt_89_to_assign_stmt_1130/slice_354_Sample/ra
      -- 
    ra_1501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_354_inst_ack_0, ack => maxPool4_CP_307_elements(278)); -- 
    -- CP-element group 279:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	277 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	357 
    -- CP-element group 279: marked-successors 
    -- CP-element group 279: 	277 
    -- CP-element group 279:  members (3) 
      -- CP-element group 279: 	 assign_stmt_89_to_assign_stmt_1130/slice_354_update_completed_
      -- CP-element group 279: 	 assign_stmt_89_to_assign_stmt_1130/slice_354_Update/$exit
      -- CP-element group 279: 	 assign_stmt_89_to_assign_stmt_1130/slice_354_Update/ca
      -- 
    ca_1506_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_354_inst_ack_1, ack => maxPool4_CP_307_elements(279)); -- 
    -- CP-element group 280:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	51 
    -- CP-element group 280: marked-predecessors 
    -- CP-element group 280: 	282 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	282 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 assign_stmt_89_to_assign_stmt_1130/slice_358_sample_start_
      -- CP-element group 280: 	 assign_stmt_89_to_assign_stmt_1130/slice_358_Sample/$entry
      -- CP-element group 280: 	 assign_stmt_89_to_assign_stmt_1130/slice_358_Sample/rr
      -- 
    rr_1514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(280), ack => slice_358_inst_req_0); -- 
    maxPool4_cp_element_group_280: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_280"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(51) & maxPool4_CP_307_elements(282);
      gj_maxPool4_cp_element_group_280 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(280), clk => clk, reset => reset); --
    end block;
    -- CP-element group 281:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: marked-predecessors 
    -- CP-element group 281: 	283 
    -- CP-element group 281: 	359 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	283 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 assign_stmt_89_to_assign_stmt_1130/slice_358_update_start_
      -- CP-element group 281: 	 assign_stmt_89_to_assign_stmt_1130/slice_358_Update/$entry
      -- CP-element group 281: 	 assign_stmt_89_to_assign_stmt_1130/slice_358_Update/cr
      -- 
    cr_1519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(281), ack => slice_358_inst_req_1); -- 
    maxPool4_cp_element_group_281: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_281"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(283) & maxPool4_CP_307_elements(359);
      gj_maxPool4_cp_element_group_281 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(281), clk => clk, reset => reset); --
    end block;
    -- CP-element group 282:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	280 
    -- CP-element group 282: successors 
    -- CP-element group 282: marked-successors 
    -- CP-element group 282: 	49 
    -- CP-element group 282: 	280 
    -- CP-element group 282:  members (3) 
      -- CP-element group 282: 	 assign_stmt_89_to_assign_stmt_1130/slice_358_sample_completed_
      -- CP-element group 282: 	 assign_stmt_89_to_assign_stmt_1130/slice_358_Sample/$exit
      -- CP-element group 282: 	 assign_stmt_89_to_assign_stmt_1130/slice_358_Sample/ra
      -- 
    ra_1515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_358_inst_ack_0, ack => maxPool4_CP_307_elements(282)); -- 
    -- CP-element group 283:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	281 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	357 
    -- CP-element group 283: marked-successors 
    -- CP-element group 283: 	281 
    -- CP-element group 283:  members (3) 
      -- CP-element group 283: 	 assign_stmt_89_to_assign_stmt_1130/slice_358_update_completed_
      -- CP-element group 283: 	 assign_stmt_89_to_assign_stmt_1130/slice_358_Update/$exit
      -- CP-element group 283: 	 assign_stmt_89_to_assign_stmt_1130/slice_358_Update/ca
      -- 
    ca_1520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 283_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_358_inst_ack_1, ack => maxPool4_CP_307_elements(283)); -- 
    -- CP-element group 284:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	51 
    -- CP-element group 284: marked-predecessors 
    -- CP-element group 284: 	286 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	286 
    -- CP-element group 284:  members (3) 
      -- CP-element group 284: 	 assign_stmt_89_to_assign_stmt_1130/slice_362_sample_start_
      -- CP-element group 284: 	 assign_stmt_89_to_assign_stmt_1130/slice_362_Sample/$entry
      -- CP-element group 284: 	 assign_stmt_89_to_assign_stmt_1130/slice_362_Sample/rr
      -- 
    rr_1528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(284), ack => slice_362_inst_req_0); -- 
    maxPool4_cp_element_group_284: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_284"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(51) & maxPool4_CP_307_elements(286);
      gj_maxPool4_cp_element_group_284 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(284), clk => clk, reset => reset); --
    end block;
    -- CP-element group 285:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: marked-predecessors 
    -- CP-element group 285: 	287 
    -- CP-element group 285: 	359 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	287 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 assign_stmt_89_to_assign_stmt_1130/slice_362_update_start_
      -- CP-element group 285: 	 assign_stmt_89_to_assign_stmt_1130/slice_362_Update/$entry
      -- CP-element group 285: 	 assign_stmt_89_to_assign_stmt_1130/slice_362_Update/cr
      -- 
    cr_1533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(285), ack => slice_362_inst_req_1); -- 
    maxPool4_cp_element_group_285: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_285"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(287) & maxPool4_CP_307_elements(359);
      gj_maxPool4_cp_element_group_285 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(285), clk => clk, reset => reset); --
    end block;
    -- CP-element group 286:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	284 
    -- CP-element group 286: successors 
    -- CP-element group 286: marked-successors 
    -- CP-element group 286: 	49 
    -- CP-element group 286: 	284 
    -- CP-element group 286:  members (3) 
      -- CP-element group 286: 	 assign_stmt_89_to_assign_stmt_1130/slice_362_sample_completed_
      -- CP-element group 286: 	 assign_stmt_89_to_assign_stmt_1130/slice_362_Sample/$exit
      -- CP-element group 286: 	 assign_stmt_89_to_assign_stmt_1130/slice_362_Sample/ra
      -- 
    ra_1529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_362_inst_ack_0, ack => maxPool4_CP_307_elements(286)); -- 
    -- CP-element group 287:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	285 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	357 
    -- CP-element group 287: marked-successors 
    -- CP-element group 287: 	285 
    -- CP-element group 287:  members (3) 
      -- CP-element group 287: 	 assign_stmt_89_to_assign_stmt_1130/slice_362_update_completed_
      -- CP-element group 287: 	 assign_stmt_89_to_assign_stmt_1130/slice_362_Update/$exit
      -- CP-element group 287: 	 assign_stmt_89_to_assign_stmt_1130/slice_362_Update/ca
      -- 
    ca_1534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_362_inst_ack_1, ack => maxPool4_CP_307_elements(287)); -- 
    -- CP-element group 288:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	51 
    -- CP-element group 288: marked-predecessors 
    -- CP-element group 288: 	290 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	290 
    -- CP-element group 288:  members (3) 
      -- CP-element group 288: 	 assign_stmt_89_to_assign_stmt_1130/slice_366_Sample/rr
      -- CP-element group 288: 	 assign_stmt_89_to_assign_stmt_1130/slice_366_Sample/$entry
      -- CP-element group 288: 	 assign_stmt_89_to_assign_stmt_1130/slice_366_sample_start_
      -- 
    rr_1542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(288), ack => slice_366_inst_req_0); -- 
    maxPool4_cp_element_group_288: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_288"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(51) & maxPool4_CP_307_elements(290);
      gj_maxPool4_cp_element_group_288 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(288), clk => clk, reset => reset); --
    end block;
    -- CP-element group 289:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: marked-predecessors 
    -- CP-element group 289: 	291 
    -- CP-element group 289: 	359 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	291 
    -- CP-element group 289:  members (3) 
      -- CP-element group 289: 	 assign_stmt_89_to_assign_stmt_1130/slice_366_Update/cr
      -- CP-element group 289: 	 assign_stmt_89_to_assign_stmt_1130/slice_366_Update/$entry
      -- CP-element group 289: 	 assign_stmt_89_to_assign_stmt_1130/slice_366_update_start_
      -- 
    cr_1547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(289), ack => slice_366_inst_req_1); -- 
    maxPool4_cp_element_group_289: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_289"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(291) & maxPool4_CP_307_elements(359);
      gj_maxPool4_cp_element_group_289 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(289), clk => clk, reset => reset); --
    end block;
    -- CP-element group 290:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	288 
    -- CP-element group 290: successors 
    -- CP-element group 290: marked-successors 
    -- CP-element group 290: 	49 
    -- CP-element group 290: 	288 
    -- CP-element group 290:  members (3) 
      -- CP-element group 290: 	 assign_stmt_89_to_assign_stmt_1130/slice_366_Sample/ra
      -- CP-element group 290: 	 assign_stmt_89_to_assign_stmt_1130/slice_366_Sample/$exit
      -- CP-element group 290: 	 assign_stmt_89_to_assign_stmt_1130/slice_366_sample_completed_
      -- 
    ra_1543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_366_inst_ack_0, ack => maxPool4_CP_307_elements(290)); -- 
    -- CP-element group 291:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	289 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	357 
    -- CP-element group 291: marked-successors 
    -- CP-element group 291: 	289 
    -- CP-element group 291:  members (3) 
      -- CP-element group 291: 	 assign_stmt_89_to_assign_stmt_1130/slice_366_Update/ca
      -- CP-element group 291: 	 assign_stmt_89_to_assign_stmt_1130/slice_366_Update/$exit
      -- CP-element group 291: 	 assign_stmt_89_to_assign_stmt_1130/slice_366_update_completed_
      -- 
    ca_1548_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_366_inst_ack_1, ack => maxPool4_CP_307_elements(291)); -- 
    -- CP-element group 292:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	51 
    -- CP-element group 292: marked-predecessors 
    -- CP-element group 292: 	294 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	294 
    -- CP-element group 292:  members (3) 
      -- CP-element group 292: 	 assign_stmt_89_to_assign_stmt_1130/slice_370_Sample/rr
      -- CP-element group 292: 	 assign_stmt_89_to_assign_stmt_1130/slice_370_Sample/$entry
      -- CP-element group 292: 	 assign_stmt_89_to_assign_stmt_1130/slice_370_sample_start_
      -- 
    rr_1556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(292), ack => slice_370_inst_req_0); -- 
    maxPool4_cp_element_group_292: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_292"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(51) & maxPool4_CP_307_elements(294);
      gj_maxPool4_cp_element_group_292 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(292), clk => clk, reset => reset); --
    end block;
    -- CP-element group 293:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: marked-predecessors 
    -- CP-element group 293: 	295 
    -- CP-element group 293: 	378 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	295 
    -- CP-element group 293:  members (3) 
      -- CP-element group 293: 	 assign_stmt_89_to_assign_stmt_1130/slice_370_Update/cr
      -- CP-element group 293: 	 assign_stmt_89_to_assign_stmt_1130/slice_370_Update/$entry
      -- CP-element group 293: 	 assign_stmt_89_to_assign_stmt_1130/slice_370_update_start_
      -- 
    cr_1561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(293), ack => slice_370_inst_req_1); -- 
    maxPool4_cp_element_group_293: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_293"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(295) & maxPool4_CP_307_elements(378);
      gj_maxPool4_cp_element_group_293 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(293), clk => clk, reset => reset); --
    end block;
    -- CP-element group 294:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	292 
    -- CP-element group 294: successors 
    -- CP-element group 294: marked-successors 
    -- CP-element group 294: 	49 
    -- CP-element group 294: 	292 
    -- CP-element group 294:  members (3) 
      -- CP-element group 294: 	 assign_stmt_89_to_assign_stmt_1130/slice_370_Sample/ra
      -- CP-element group 294: 	 assign_stmt_89_to_assign_stmt_1130/slice_370_Sample/$exit
      -- CP-element group 294: 	 assign_stmt_89_to_assign_stmt_1130/slice_370_sample_completed_
      -- 
    ra_1557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 294_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_370_inst_ack_0, ack => maxPool4_CP_307_elements(294)); -- 
    -- CP-element group 295:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	293 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	376 
    -- CP-element group 295: marked-successors 
    -- CP-element group 295: 	293 
    -- CP-element group 295:  members (3) 
      -- CP-element group 295: 	 assign_stmt_89_to_assign_stmt_1130/slice_370_Update/ca
      -- CP-element group 295: 	 assign_stmt_89_to_assign_stmt_1130/slice_370_Update/$exit
      -- CP-element group 295: 	 assign_stmt_89_to_assign_stmt_1130/slice_370_update_completed_
      -- 
    ca_1562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_370_inst_ack_1, ack => maxPool4_CP_307_elements(295)); -- 
    -- CP-element group 296:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	51 
    -- CP-element group 296: marked-predecessors 
    -- CP-element group 296: 	298 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	298 
    -- CP-element group 296:  members (3) 
      -- CP-element group 296: 	 assign_stmt_89_to_assign_stmt_1130/slice_374_Sample/rr
      -- CP-element group 296: 	 assign_stmt_89_to_assign_stmt_1130/slice_374_Sample/$entry
      -- CP-element group 296: 	 assign_stmt_89_to_assign_stmt_1130/slice_374_sample_start_
      -- 
    rr_1570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(296), ack => slice_374_inst_req_0); -- 
    maxPool4_cp_element_group_296: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_296"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(51) & maxPool4_CP_307_elements(298);
      gj_maxPool4_cp_element_group_296 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(296), clk => clk, reset => reset); --
    end block;
    -- CP-element group 297:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: marked-predecessors 
    -- CP-element group 297: 	299 
    -- CP-element group 297: 	378 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	299 
    -- CP-element group 297:  members (3) 
      -- CP-element group 297: 	 assign_stmt_89_to_assign_stmt_1130/slice_374_Update/$entry
      -- CP-element group 297: 	 assign_stmt_89_to_assign_stmt_1130/slice_374_Update/cr
      -- CP-element group 297: 	 assign_stmt_89_to_assign_stmt_1130/slice_374_update_start_
      -- 
    cr_1575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(297), ack => slice_374_inst_req_1); -- 
    maxPool4_cp_element_group_297: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_297"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(299) & maxPool4_CP_307_elements(378);
      gj_maxPool4_cp_element_group_297 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(297), clk => clk, reset => reset); --
    end block;
    -- CP-element group 298:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	296 
    -- CP-element group 298: successors 
    -- CP-element group 298: marked-successors 
    -- CP-element group 298: 	49 
    -- CP-element group 298: 	296 
    -- CP-element group 298:  members (3) 
      -- CP-element group 298: 	 assign_stmt_89_to_assign_stmt_1130/slice_374_Sample/ra
      -- CP-element group 298: 	 assign_stmt_89_to_assign_stmt_1130/slice_374_Sample/$exit
      -- CP-element group 298: 	 assign_stmt_89_to_assign_stmt_1130/slice_374_sample_completed_
      -- 
    ra_1571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 298_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_374_inst_ack_0, ack => maxPool4_CP_307_elements(298)); -- 
    -- CP-element group 299:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	297 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	376 
    -- CP-element group 299: marked-successors 
    -- CP-element group 299: 	297 
    -- CP-element group 299:  members (3) 
      -- CP-element group 299: 	 assign_stmt_89_to_assign_stmt_1130/slice_374_Update/ca
      -- CP-element group 299: 	 assign_stmt_89_to_assign_stmt_1130/slice_374_Update/$exit
      -- CP-element group 299: 	 assign_stmt_89_to_assign_stmt_1130/slice_374_update_completed_
      -- 
    ca_1576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_374_inst_ack_1, ack => maxPool4_CP_307_elements(299)); -- 
    -- CP-element group 300:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	51 
    -- CP-element group 300: marked-predecessors 
    -- CP-element group 300: 	302 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	302 
    -- CP-element group 300:  members (3) 
      -- CP-element group 300: 	 assign_stmt_89_to_assign_stmt_1130/slice_378_sample_start_
      -- CP-element group 300: 	 assign_stmt_89_to_assign_stmt_1130/slice_378_Sample/$entry
      -- CP-element group 300: 	 assign_stmt_89_to_assign_stmt_1130/slice_378_Sample/rr
      -- 
    rr_1584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(300), ack => slice_378_inst_req_0); -- 
    maxPool4_cp_element_group_300: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_300"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(51) & maxPool4_CP_307_elements(302);
      gj_maxPool4_cp_element_group_300 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(300), clk => clk, reset => reset); --
    end block;
    -- CP-element group 301:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: marked-predecessors 
    -- CP-element group 301: 	303 
    -- CP-element group 301: 	378 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	303 
    -- CP-element group 301:  members (3) 
      -- CP-element group 301: 	 assign_stmt_89_to_assign_stmt_1130/slice_378_update_start_
      -- CP-element group 301: 	 assign_stmt_89_to_assign_stmt_1130/slice_378_Update/$entry
      -- CP-element group 301: 	 assign_stmt_89_to_assign_stmt_1130/slice_378_Update/cr
      -- 
    cr_1589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(301), ack => slice_378_inst_req_1); -- 
    maxPool4_cp_element_group_301: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_301"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(303) & maxPool4_CP_307_elements(378);
      gj_maxPool4_cp_element_group_301 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(301), clk => clk, reset => reset); --
    end block;
    -- CP-element group 302:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	300 
    -- CP-element group 302: successors 
    -- CP-element group 302: marked-successors 
    -- CP-element group 302: 	49 
    -- CP-element group 302: 	300 
    -- CP-element group 302:  members (3) 
      -- CP-element group 302: 	 assign_stmt_89_to_assign_stmt_1130/slice_378_sample_completed_
      -- CP-element group 302: 	 assign_stmt_89_to_assign_stmt_1130/slice_378_Sample/$exit
      -- CP-element group 302: 	 assign_stmt_89_to_assign_stmt_1130/slice_378_Sample/ra
      -- 
    ra_1585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 302_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_378_inst_ack_0, ack => maxPool4_CP_307_elements(302)); -- 
    -- CP-element group 303:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	301 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	376 
    -- CP-element group 303: marked-successors 
    -- CP-element group 303: 	301 
    -- CP-element group 303:  members (3) 
      -- CP-element group 303: 	 assign_stmt_89_to_assign_stmt_1130/slice_378_update_completed_
      -- CP-element group 303: 	 assign_stmt_89_to_assign_stmt_1130/slice_378_Update/$exit
      -- CP-element group 303: 	 assign_stmt_89_to_assign_stmt_1130/slice_378_Update/ca
      -- 
    ca_1590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_378_inst_ack_1, ack => maxPool4_CP_307_elements(303)); -- 
    -- CP-element group 304:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	51 
    -- CP-element group 304: marked-predecessors 
    -- CP-element group 304: 	306 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	306 
    -- CP-element group 304:  members (3) 
      -- CP-element group 304: 	 assign_stmt_89_to_assign_stmt_1130/slice_382_sample_start_
      -- CP-element group 304: 	 assign_stmt_89_to_assign_stmt_1130/slice_382_Sample/$entry
      -- CP-element group 304: 	 assign_stmt_89_to_assign_stmt_1130/slice_382_Sample/rr
      -- 
    rr_1598_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1598_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(304), ack => slice_382_inst_req_0); -- 
    maxPool4_cp_element_group_304: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_304"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(51) & maxPool4_CP_307_elements(306);
      gj_maxPool4_cp_element_group_304 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(304), clk => clk, reset => reset); --
    end block;
    -- CP-element group 305:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: marked-predecessors 
    -- CP-element group 305: 	307 
    -- CP-element group 305: 	378 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	307 
    -- CP-element group 305:  members (3) 
      -- CP-element group 305: 	 assign_stmt_89_to_assign_stmt_1130/slice_382_Update/cr
      -- CP-element group 305: 	 assign_stmt_89_to_assign_stmt_1130/slice_382_update_start_
      -- CP-element group 305: 	 assign_stmt_89_to_assign_stmt_1130/slice_382_Update/$entry
      -- 
    cr_1603_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1603_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(305), ack => slice_382_inst_req_1); -- 
    maxPool4_cp_element_group_305: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_305"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(307) & maxPool4_CP_307_elements(378);
      gj_maxPool4_cp_element_group_305 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(305), clk => clk, reset => reset); --
    end block;
    -- CP-element group 306:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	304 
    -- CP-element group 306: successors 
    -- CP-element group 306: marked-successors 
    -- CP-element group 306: 	49 
    -- CP-element group 306: 	304 
    -- CP-element group 306:  members (3) 
      -- CP-element group 306: 	 assign_stmt_89_to_assign_stmt_1130/slice_382_sample_completed_
      -- CP-element group 306: 	 assign_stmt_89_to_assign_stmt_1130/slice_382_Sample/$exit
      -- CP-element group 306: 	 assign_stmt_89_to_assign_stmt_1130/slice_382_Sample/ra
      -- 
    ra_1599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_382_inst_ack_0, ack => maxPool4_CP_307_elements(306)); -- 
    -- CP-element group 307:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	305 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	376 
    -- CP-element group 307: marked-successors 
    -- CP-element group 307: 	305 
    -- CP-element group 307:  members (3) 
      -- CP-element group 307: 	 assign_stmt_89_to_assign_stmt_1130/slice_382_Update/$exit
      -- CP-element group 307: 	 assign_stmt_89_to_assign_stmt_1130/slice_382_Update/ca
      -- CP-element group 307: 	 assign_stmt_89_to_assign_stmt_1130/slice_382_update_completed_
      -- 
    ca_1604_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_382_inst_ack_1, ack => maxPool4_CP_307_elements(307)); -- 
    -- CP-element group 308:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	312 
    -- CP-element group 308: marked-predecessors 
    -- CP-element group 308: 	313 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	313 
    -- CP-element group 308:  members (3) 
      -- CP-element group 308: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1030_request/req
      -- CP-element group 308: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1030_sample_start_
      -- CP-element group 308: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1030_request/$entry
      -- 
    req_1644_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1644_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(308), ack => addr_of_1030_final_reg_req_0); -- 
    maxPool4_cp_element_group_308: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_308"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(312) & maxPool4_CP_307_elements(313);
      gj_maxPool4_cp_element_group_308 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(308), clk => clk, reset => reset); --
    end block;
    -- CP-element group 309:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	1 
    -- CP-element group 309: marked-predecessors 
    -- CP-element group 309: 	314 
    -- CP-element group 309: 	317 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	314 
    -- CP-element group 309:  members (3) 
      -- CP-element group 309: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1030_update_start_
      -- CP-element group 309: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1030_complete/$entry
      -- CP-element group 309: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1030_complete/req
      -- 
    req_1649_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1649_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(309), ack => addr_of_1030_final_reg_req_1); -- 
    maxPool4_cp_element_group_309: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_309"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(1) & maxPool4_CP_307_elements(314) & maxPool4_CP_307_elements(317);
      gj_maxPool4_cp_element_group_309 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(309), clk => clk, reset => reset); --
    end block;
    -- CP-element group 310:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	1 
    -- CP-element group 310: marked-predecessors 
    -- CP-element group 310: 	312 
    -- CP-element group 310: 	313 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	312 
    -- CP-element group 310:  members (3) 
      -- CP-element group 310: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1029_final_index_sum_regn_Update/req
      -- CP-element group 310: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1029_final_index_sum_regn_Update/$entry
      -- CP-element group 310: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1029_final_index_sum_regn_update_start
      -- 
    req_1634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(310), ack => array_obj_ref_1029_index_offset_req_1); -- 
    maxPool4_cp_element_group_310: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_310"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(1) & maxPool4_CP_307_elements(312) & maxPool4_CP_307_elements(313);
      gj_maxPool4_cp_element_group_310 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(310), clk => clk, reset => reset); --
    end block;
    -- CP-element group 311:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	1 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	391 
    -- CP-element group 311: marked-successors 
    -- CP-element group 311: 	2 
    -- CP-element group 311:  members (3) 
      -- CP-element group 311: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1029_final_index_sum_regn_Sample/ack
      -- CP-element group 311: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1029_final_index_sum_regn_Sample/$exit
      -- CP-element group 311: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1029_final_index_sum_regn_sample_complete
      -- 
    ack_1630_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1029_index_offset_ack_0, ack => maxPool4_CP_307_elements(311)); -- 
    -- CP-element group 312:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	310 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	308 
    -- CP-element group 312: marked-successors 
    -- CP-element group 312: 	310 
    -- CP-element group 312:  members (8) 
      -- CP-element group 312: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1029_offset_calculated
      -- CP-element group 312: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1029_root_address_calculated
      -- CP-element group 312: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1029_base_plus_offset/sum_rename_ack
      -- CP-element group 312: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1029_base_plus_offset/sum_rename_req
      -- CP-element group 312: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1029_base_plus_offset/$exit
      -- CP-element group 312: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1029_base_plus_offset/$entry
      -- CP-element group 312: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1029_final_index_sum_regn_Update/ack
      -- CP-element group 312: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1029_final_index_sum_regn_Update/$exit
      -- 
    ack_1635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1029_index_offset_ack_1, ack => maxPool4_CP_307_elements(312)); -- 
    -- CP-element group 313:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	308 
    -- CP-element group 313: successors 
    -- CP-element group 313: marked-successors 
    -- CP-element group 313: 	308 
    -- CP-element group 313: 	310 
    -- CP-element group 313:  members (3) 
      -- CP-element group 313: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1030_sample_completed_
      -- CP-element group 313: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1030_request/ack
      -- CP-element group 313: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1030_request/$exit
      -- 
    ack_1645_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1030_final_reg_ack_0, ack => maxPool4_CP_307_elements(313)); -- 
    -- CP-element group 314:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	309 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	315 
    -- CP-element group 314: marked-successors 
    -- CP-element group 314: 	309 
    -- CP-element group 314:  members (3) 
      -- CP-element group 314: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1030_complete/$exit
      -- CP-element group 314: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1030_complete/ack
      -- CP-element group 314: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1030_update_completed_
      -- 
    ack_1650_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1030_final_reg_ack_1, ack => maxPool4_CP_307_elements(314)); -- 
    -- CP-element group 315:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	314 
    -- CP-element group 315: marked-predecessors 
    -- CP-element group 315: 	317 
    -- CP-element group 315: successors 
    -- CP-element group 315: 	317 
    -- CP-element group 315:  members (3) 
      -- CP-element group 315: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1034_sample_start_
      -- CP-element group 315: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1034_Sample/$entry
      -- CP-element group 315: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1034_Sample/req
      -- 
    req_1658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(315), ack => W_myptr5_1032_delayed_8_0_1032_inst_req_0); -- 
    maxPool4_cp_element_group_315: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_315"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(314) & maxPool4_CP_307_elements(317);
      gj_maxPool4_cp_element_group_315 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(315), clk => clk, reset => reset); --
    end block;
    -- CP-element group 316:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: marked-predecessors 
    -- CP-element group 316: 	318 
    -- CP-element group 316: 	325 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	318 
    -- CP-element group 316:  members (3) 
      -- CP-element group 316: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1034_update_start_
      -- CP-element group 316: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1034_Update/$entry
      -- CP-element group 316: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1034_Update/req
      -- 
    req_1663_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1663_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(316), ack => W_myptr5_1032_delayed_8_0_1032_inst_req_1); -- 
    maxPool4_cp_element_group_316: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_316"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(318) & maxPool4_CP_307_elements(325);
      gj_maxPool4_cp_element_group_316 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(316), clk => clk, reset => reset); --
    end block;
    -- CP-element group 317:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	315 
    -- CP-element group 317: successors 
    -- CP-element group 317: marked-successors 
    -- CP-element group 317: 	309 
    -- CP-element group 317: 	315 
    -- CP-element group 317:  members (3) 
      -- CP-element group 317: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1034_sample_completed_
      -- CP-element group 317: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1034_Sample/$exit
      -- CP-element group 317: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1034_Sample/ack
      -- 
    ack_1659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 317_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_myptr5_1032_delayed_8_0_1032_inst_ack_0, ack => maxPool4_CP_307_elements(317)); -- 
    -- CP-element group 318:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	316 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	323 
    -- CP-element group 318: marked-successors 
    -- CP-element group 318: 	316 
    -- CP-element group 318:  members (19) 
      -- CP-element group 318: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1036_base_address_calculated
      -- CP-element group 318: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1036_word_address_calculated
      -- CP-element group 318: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1036_root_address_calculated
      -- CP-element group 318: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1036_base_plus_offset/sum_rename_req
      -- CP-element group 318: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1036_base_plus_offset/sum_rename_ack
      -- CP-element group 318: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1036_word_addrgen/$entry
      -- CP-element group 318: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1036_word_addrgen/$exit
      -- CP-element group 318: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1036_base_address_resized
      -- CP-element group 318: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1036_base_addr_resize/$entry
      -- CP-element group 318: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1034_update_completed_
      -- CP-element group 318: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1034_Update/$exit
      -- CP-element group 318: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1034_Update/ack
      -- CP-element group 318: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1036_base_addr_resize/$exit
      -- CP-element group 318: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1036_base_addr_resize/base_resize_req
      -- CP-element group 318: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1036_base_addr_resize/base_resize_ack
      -- CP-element group 318: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1036_base_plus_offset/$entry
      -- CP-element group 318: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1036_base_plus_offset/$exit
      -- CP-element group 318: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1036_word_addrgen/root_register_req
      -- CP-element group 318: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1036_word_addrgen/root_register_ack
      -- 
    ack_1664_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 318_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_myptr5_1032_delayed_8_0_1032_inst_ack_1, ack => maxPool4_CP_307_elements(318)); -- 
    -- CP-element group 319:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	55 
    -- CP-element group 319: 	59 
    -- CP-element group 319: 	63 
    -- CP-element group 319: 	67 
    -- CP-element group 319: 	119 
    -- CP-element group 319: 	123 
    -- CP-element group 319: 	127 
    -- CP-element group 319: 	131 
    -- CP-element group 319: 	183 
    -- CP-element group 319: 	187 
    -- CP-element group 319: 	191 
    -- CP-element group 319: 	195 
    -- CP-element group 319: 	247 
    -- CP-element group 319: 	251 
    -- CP-element group 319: 	255 
    -- CP-element group 319: 	259 
    -- CP-element group 319: marked-predecessors 
    -- CP-element group 319: 	321 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	321 
    -- CP-element group 319:  members (3) 
      -- CP-element group 319: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1047_sample_start_
      -- CP-element group 319: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1047_Sample/$entry
      -- CP-element group 319: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1047_Sample/rr
      -- 
    rr_1672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(319), ack => CONCAT_u32_u64_1047_inst_req_0); -- 
    maxPool4_cp_element_group_319: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 1);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_319"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(55) & maxPool4_CP_307_elements(59) & maxPool4_CP_307_elements(63) & maxPool4_CP_307_elements(67) & maxPool4_CP_307_elements(119) & maxPool4_CP_307_elements(123) & maxPool4_CP_307_elements(127) & maxPool4_CP_307_elements(131) & maxPool4_CP_307_elements(183) & maxPool4_CP_307_elements(187) & maxPool4_CP_307_elements(191) & maxPool4_CP_307_elements(195) & maxPool4_CP_307_elements(247) & maxPool4_CP_307_elements(251) & maxPool4_CP_307_elements(255) & maxPool4_CP_307_elements(259) & maxPool4_CP_307_elements(321);
      gj_maxPool4_cp_element_group_319 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(319), clk => clk, reset => reset); --
    end block;
    -- CP-element group 320:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: marked-predecessors 
    -- CP-element group 320: 	322 
    -- CP-element group 320: 	325 
    -- CP-element group 320: successors 
    -- CP-element group 320: 	322 
    -- CP-element group 320:  members (3) 
      -- CP-element group 320: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1047_update_start_
      -- CP-element group 320: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1047_Update/$entry
      -- CP-element group 320: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1047_Update/cr
      -- 
    cr_1677_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1677_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(320), ack => CONCAT_u32_u64_1047_inst_req_1); -- 
    maxPool4_cp_element_group_320: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_320"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(322) & maxPool4_CP_307_elements(325);
      gj_maxPool4_cp_element_group_320 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(320), clk => clk, reset => reset); --
    end block;
    -- CP-element group 321:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	319 
    -- CP-element group 321: successors 
    -- CP-element group 321: marked-successors 
    -- CP-element group 321: 	53 
    -- CP-element group 321: 	57 
    -- CP-element group 321: 	61 
    -- CP-element group 321: 	65 
    -- CP-element group 321: 	117 
    -- CP-element group 321: 	121 
    -- CP-element group 321: 	125 
    -- CP-element group 321: 	129 
    -- CP-element group 321: 	181 
    -- CP-element group 321: 	185 
    -- CP-element group 321: 	189 
    -- CP-element group 321: 	193 
    -- CP-element group 321: 	245 
    -- CP-element group 321: 	249 
    -- CP-element group 321: 	253 
    -- CP-element group 321: 	257 
    -- CP-element group 321: 	319 
    -- CP-element group 321:  members (3) 
      -- CP-element group 321: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1047_sample_completed_
      -- CP-element group 321: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1047_Sample/$exit
      -- CP-element group 321: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1047_Sample/ra
      -- 
    ra_1673_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_1047_inst_ack_0, ack => maxPool4_CP_307_elements(321)); -- 
    -- CP-element group 322:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	320 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	323 
    -- CP-element group 322: marked-successors 
    -- CP-element group 322: 	320 
    -- CP-element group 322:  members (3) 
      -- CP-element group 322: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1047_Update/ca
      -- CP-element group 322: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1047_update_completed_
      -- CP-element group 322: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1047_Update/$exit
      -- 
    ca_1678_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 322_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_1047_inst_ack_1, ack => maxPool4_CP_307_elements(322)); -- 
    -- CP-element group 323:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	318 
    -- CP-element group 323: 	322 
    -- CP-element group 323: marked-predecessors 
    -- CP-element group 323: 	325 
    -- CP-element group 323: 	382 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	325 
    -- CP-element group 323:  members (9) 
      -- CP-element group 323: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1036_Sample/word_access_start/word_0/$entry
      -- CP-element group 323: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1036_sample_start_
      -- CP-element group 323: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1036_Sample/word_access_start/word_0/rr
      -- CP-element group 323: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1036_Sample/$entry
      -- CP-element group 323: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1036_Sample/word_access_start/$entry
      -- CP-element group 323: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1036_Sample/ptr_deref_1036_Split/$entry
      -- CP-element group 323: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1036_Sample/ptr_deref_1036_Split/$exit
      -- CP-element group 323: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1036_Sample/ptr_deref_1036_Split/split_req
      -- CP-element group 323: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1036_Sample/ptr_deref_1036_Split/split_ack
      -- 
    rr_1716_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1716_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(323), ack => ptr_deref_1036_store_0_req_0); -- 
    maxPool4_cp_element_group_323: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_323"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(318) & maxPool4_CP_307_elements(322) & maxPool4_CP_307_elements(325) & maxPool4_CP_307_elements(382);
      gj_maxPool4_cp_element_group_323 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(323), clk => clk, reset => reset); --
    end block;
    -- CP-element group 324:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: marked-predecessors 
    -- CP-element group 324: 	326 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	326 
    -- CP-element group 324:  members (5) 
      -- CP-element group 324: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1036_Update/$entry
      -- CP-element group 324: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1036_Update/word_access_complete/word_0/cr
      -- CP-element group 324: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1036_Update/word_access_complete/$entry
      -- CP-element group 324: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1036_update_start_
      -- CP-element group 324: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1036_Update/word_access_complete/word_0/$entry
      -- 
    cr_1727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(324), ack => ptr_deref_1036_store_0_req_1); -- 
    maxPool4_cp_element_group_324: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_324"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_307_elements(326);
      gj_maxPool4_cp_element_group_324 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(324), clk => clk, reset => reset); --
    end block;
    -- CP-element group 325:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	323 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	388 
    -- CP-element group 325: marked-successors 
    -- CP-element group 325: 	316 
    -- CP-element group 325: 	320 
    -- CP-element group 325: 	323 
    -- CP-element group 325:  members (5) 
      -- CP-element group 325: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1036_Sample/word_access_start/word_0/ra
      -- CP-element group 325: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1036_sample_completed_
      -- CP-element group 325: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1036_Sample/word_access_start/word_0/$exit
      -- CP-element group 325: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1036_Sample/word_access_start/$exit
      -- CP-element group 325: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1036_Sample/$exit
      -- 
    ra_1717_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 325_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1036_store_0_ack_0, ack => maxPool4_CP_307_elements(325)); -- 
    -- CP-element group 326:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	324 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	391 
    -- CP-element group 326: marked-successors 
    -- CP-element group 326: 	324 
    -- CP-element group 326:  members (5) 
      -- CP-element group 326: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1036_Update/word_access_complete/word_0/$exit
      -- CP-element group 326: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1036_update_completed_
      -- CP-element group 326: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1036_Update/$exit
      -- CP-element group 326: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1036_Update/word_access_complete/word_0/ca
      -- CP-element group 326: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1036_Update/word_access_complete/$exit
      -- 
    ca_1728_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 326_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1036_store_0_ack_1, ack => maxPool4_CP_307_elements(326)); -- 
    -- CP-element group 327:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	331 
    -- CP-element group 327: marked-predecessors 
    -- CP-element group 327: 	332 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	332 
    -- CP-element group 327:  members (3) 
      -- CP-element group 327: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1056_sample_start_
      -- CP-element group 327: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1056_request/req
      -- CP-element group 327: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1056_request/$entry
      -- 
    req_1768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(327), ack => addr_of_1056_final_reg_req_0); -- 
    maxPool4_cp_element_group_327: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_327"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(331) & maxPool4_CP_307_elements(332);
      gj_maxPool4_cp_element_group_327 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(327), clk => clk, reset => reset); --
    end block;
    -- CP-element group 328:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	1 
    -- CP-element group 328: marked-predecessors 
    -- CP-element group 328: 	333 
    -- CP-element group 328: 	336 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	333 
    -- CP-element group 328:  members (3) 
      -- CP-element group 328: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1056_update_start_
      -- CP-element group 328: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1056_complete/req
      -- CP-element group 328: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1056_complete/$entry
      -- 
    req_1773_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1773_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(328), ack => addr_of_1056_final_reg_req_1); -- 
    maxPool4_cp_element_group_328: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_328"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(1) & maxPool4_CP_307_elements(333) & maxPool4_CP_307_elements(336);
      gj_maxPool4_cp_element_group_328 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(328), clk => clk, reset => reset); --
    end block;
    -- CP-element group 329:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	1 
    -- CP-element group 329: marked-predecessors 
    -- CP-element group 329: 	331 
    -- CP-element group 329: 	332 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	331 
    -- CP-element group 329:  members (3) 
      -- CP-element group 329: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1055_final_index_sum_regn_update_start
      -- CP-element group 329: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1055_final_index_sum_regn_Update/$entry
      -- CP-element group 329: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1055_final_index_sum_regn_Update/req
      -- 
    req_1758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(329), ack => array_obj_ref_1055_index_offset_req_1); -- 
    maxPool4_cp_element_group_329: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_329"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(1) & maxPool4_CP_307_elements(331) & maxPool4_CP_307_elements(332);
      gj_maxPool4_cp_element_group_329 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(329), clk => clk, reset => reset); --
    end block;
    -- CP-element group 330:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	1 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	391 
    -- CP-element group 330: marked-successors 
    -- CP-element group 330: 	2 
    -- CP-element group 330:  members (3) 
      -- CP-element group 330: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1055_final_index_sum_regn_Sample/$exit
      -- CP-element group 330: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1055_final_index_sum_regn_sample_complete
      -- CP-element group 330: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1055_final_index_sum_regn_Sample/ack
      -- 
    ack_1754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 330_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1055_index_offset_ack_0, ack => maxPool4_CP_307_elements(330)); -- 
    -- CP-element group 331:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	329 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	327 
    -- CP-element group 331: marked-successors 
    -- CP-element group 331: 	329 
    -- CP-element group 331:  members (8) 
      -- CP-element group 331: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1055_base_plus_offset/sum_rename_ack
      -- CP-element group 331: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1055_root_address_calculated
      -- CP-element group 331: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1055_offset_calculated
      -- CP-element group 331: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1055_final_index_sum_regn_Update/$exit
      -- CP-element group 331: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1055_final_index_sum_regn_Update/ack
      -- CP-element group 331: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1055_base_plus_offset/$entry
      -- CP-element group 331: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1055_base_plus_offset/$exit
      -- CP-element group 331: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1055_base_plus_offset/sum_rename_req
      -- 
    ack_1759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 331_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1055_index_offset_ack_1, ack => maxPool4_CP_307_elements(331)); -- 
    -- CP-element group 332:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	327 
    -- CP-element group 332: successors 
    -- CP-element group 332: marked-successors 
    -- CP-element group 332: 	327 
    -- CP-element group 332: 	329 
    -- CP-element group 332:  members (3) 
      -- CP-element group 332: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1056_sample_completed_
      -- CP-element group 332: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1056_request/ack
      -- CP-element group 332: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1056_request/$exit
      -- 
    ack_1769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1056_final_reg_ack_0, ack => maxPool4_CP_307_elements(332)); -- 
    -- CP-element group 333:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	328 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	334 
    -- CP-element group 333: marked-successors 
    -- CP-element group 333: 	328 
    -- CP-element group 333:  members (3) 
      -- CP-element group 333: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1056_update_completed_
      -- CP-element group 333: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1056_complete/ack
      -- CP-element group 333: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1056_complete/$exit
      -- 
    ack_1774_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 333_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1056_final_reg_ack_1, ack => maxPool4_CP_307_elements(333)); -- 
    -- CP-element group 334:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	333 
    -- CP-element group 334: marked-predecessors 
    -- CP-element group 334: 	336 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	336 
    -- CP-element group 334:  members (3) 
      -- CP-element group 334: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1060_sample_start_
      -- CP-element group 334: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1060_Sample/$entry
      -- CP-element group 334: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1060_Sample/req
      -- 
    req_1782_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1782_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(334), ack => W_myptr6_1055_delayed_8_0_1058_inst_req_0); -- 
    maxPool4_cp_element_group_334: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_334"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(333) & maxPool4_CP_307_elements(336);
      gj_maxPool4_cp_element_group_334 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(334), clk => clk, reset => reset); --
    end block;
    -- CP-element group 335:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: marked-predecessors 
    -- CP-element group 335: 	337 
    -- CP-element group 335: 	344 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	337 
    -- CP-element group 335:  members (3) 
      -- CP-element group 335: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1060_Update/req
      -- CP-element group 335: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1060_update_start_
      -- CP-element group 335: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1060_Update/$entry
      -- 
    req_1787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(335), ack => W_myptr6_1055_delayed_8_0_1058_inst_req_1); -- 
    maxPool4_cp_element_group_335: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_335"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(337) & maxPool4_CP_307_elements(344);
      gj_maxPool4_cp_element_group_335 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(335), clk => clk, reset => reset); --
    end block;
    -- CP-element group 336:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	334 
    -- CP-element group 336: successors 
    -- CP-element group 336: marked-successors 
    -- CP-element group 336: 	328 
    -- CP-element group 336: 	334 
    -- CP-element group 336:  members (3) 
      -- CP-element group 336: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1060_sample_completed_
      -- CP-element group 336: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1060_Sample/$exit
      -- CP-element group 336: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1060_Sample/ack
      -- 
    ack_1783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_myptr6_1055_delayed_8_0_1058_inst_ack_0, ack => maxPool4_CP_307_elements(336)); -- 
    -- CP-element group 337:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	335 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	342 
    -- CP-element group 337: marked-successors 
    -- CP-element group 337: 	335 
    -- CP-element group 337:  members (19) 
      -- CP-element group 337: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1062_word_addrgen/$entry
      -- CP-element group 337: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1062_word_addrgen/$exit
      -- CP-element group 337: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1060_update_completed_
      -- CP-element group 337: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1062_word_addrgen/root_register_req
      -- CP-element group 337: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1062_word_addrgen/root_register_ack
      -- CP-element group 337: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1060_Update/$exit
      -- CP-element group 337: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1062_base_address_calculated
      -- CP-element group 337: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1062_base_plus_offset/sum_rename_ack
      -- CP-element group 337: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1062_base_plus_offset/sum_rename_req
      -- CP-element group 337: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1062_base_plus_offset/$exit
      -- CP-element group 337: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1062_base_plus_offset/$entry
      -- CP-element group 337: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1062_base_addr_resize/base_resize_ack
      -- CP-element group 337: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1062_base_addr_resize/base_resize_req
      -- CP-element group 337: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1062_base_addr_resize/$exit
      -- CP-element group 337: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1062_base_addr_resize/$entry
      -- CP-element group 337: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1062_base_address_resized
      -- CP-element group 337: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1062_root_address_calculated
      -- CP-element group 337: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1060_Update/ack
      -- CP-element group 337: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1062_word_address_calculated
      -- 
    ack_1788_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_myptr6_1055_delayed_8_0_1058_inst_ack_1, ack => maxPool4_CP_307_elements(337)); -- 
    -- CP-element group 338:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	71 
    -- CP-element group 338: 	75 
    -- CP-element group 338: 	79 
    -- CP-element group 338: 	83 
    -- CP-element group 338: 	135 
    -- CP-element group 338: 	139 
    -- CP-element group 338: 	143 
    -- CP-element group 338: 	147 
    -- CP-element group 338: 	199 
    -- CP-element group 338: 	203 
    -- CP-element group 338: 	207 
    -- CP-element group 338: 	211 
    -- CP-element group 338: 	263 
    -- CP-element group 338: 	267 
    -- CP-element group 338: 	271 
    -- CP-element group 338: 	275 
    -- CP-element group 338: marked-predecessors 
    -- CP-element group 338: 	340 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	340 
    -- CP-element group 338:  members (3) 
      -- CP-element group 338: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1073_Sample/$entry
      -- CP-element group 338: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1073_sample_start_
      -- CP-element group 338: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1073_Sample/rr
      -- 
    rr_1796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(338), ack => CONCAT_u32_u64_1073_inst_req_0); -- 
    maxPool4_cp_element_group_338: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 1);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_338"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(71) & maxPool4_CP_307_elements(75) & maxPool4_CP_307_elements(79) & maxPool4_CP_307_elements(83) & maxPool4_CP_307_elements(135) & maxPool4_CP_307_elements(139) & maxPool4_CP_307_elements(143) & maxPool4_CP_307_elements(147) & maxPool4_CP_307_elements(199) & maxPool4_CP_307_elements(203) & maxPool4_CP_307_elements(207) & maxPool4_CP_307_elements(211) & maxPool4_CP_307_elements(263) & maxPool4_CP_307_elements(267) & maxPool4_CP_307_elements(271) & maxPool4_CP_307_elements(275) & maxPool4_CP_307_elements(340);
      gj_maxPool4_cp_element_group_338 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(338), clk => clk, reset => reset); --
    end block;
    -- CP-element group 339:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: marked-predecessors 
    -- CP-element group 339: 	341 
    -- CP-element group 339: 	344 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	341 
    -- CP-element group 339:  members (3) 
      -- CP-element group 339: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1073_Update/cr
      -- CP-element group 339: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1073_Update/$entry
      -- CP-element group 339: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1073_update_start_
      -- 
    cr_1801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(339), ack => CONCAT_u32_u64_1073_inst_req_1); -- 
    maxPool4_cp_element_group_339: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_339"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(341) & maxPool4_CP_307_elements(344);
      gj_maxPool4_cp_element_group_339 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(339), clk => clk, reset => reset); --
    end block;
    -- CP-element group 340:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	338 
    -- CP-element group 340: successors 
    -- CP-element group 340: marked-successors 
    -- CP-element group 340: 	69 
    -- CP-element group 340: 	73 
    -- CP-element group 340: 	77 
    -- CP-element group 340: 	81 
    -- CP-element group 340: 	133 
    -- CP-element group 340: 	137 
    -- CP-element group 340: 	141 
    -- CP-element group 340: 	145 
    -- CP-element group 340: 	197 
    -- CP-element group 340: 	201 
    -- CP-element group 340: 	205 
    -- CP-element group 340: 	209 
    -- CP-element group 340: 	261 
    -- CP-element group 340: 	265 
    -- CP-element group 340: 	269 
    -- CP-element group 340: 	273 
    -- CP-element group 340: 	338 
    -- CP-element group 340:  members (3) 
      -- CP-element group 340: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1073_Sample/$exit
      -- CP-element group 340: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1073_sample_completed_
      -- CP-element group 340: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1073_Sample/ra
      -- 
    ra_1797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_1073_inst_ack_0, ack => maxPool4_CP_307_elements(340)); -- 
    -- CP-element group 341:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	339 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	342 
    -- CP-element group 341: marked-successors 
    -- CP-element group 341: 	339 
    -- CP-element group 341:  members (3) 
      -- CP-element group 341: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1073_Update/$exit
      -- CP-element group 341: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1073_Update/ca
      -- CP-element group 341: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1073_update_completed_
      -- 
    ca_1802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_1073_inst_ack_1, ack => maxPool4_CP_307_elements(341)); -- 
    -- CP-element group 342:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	337 
    -- CP-element group 342: 	341 
    -- CP-element group 342: 	388 
    -- CP-element group 342: marked-predecessors 
    -- CP-element group 342: 	344 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	344 
    -- CP-element group 342:  members (9) 
      -- CP-element group 342: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1062_Sample/ptr_deref_1062_Split/$entry
      -- CP-element group 342: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1062_Sample/word_access_start/word_0/rr
      -- CP-element group 342: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1062_Sample/ptr_deref_1062_Split/$exit
      -- CP-element group 342: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1062_Sample/word_access_start/word_0/$entry
      -- CP-element group 342: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1062_sample_start_
      -- CP-element group 342: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1062_Sample/$entry
      -- CP-element group 342: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1062_Sample/ptr_deref_1062_Split/split_req
      -- CP-element group 342: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1062_Sample/ptr_deref_1062_Split/split_ack
      -- CP-element group 342: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1062_Sample/word_access_start/$entry
      -- 
    rr_1840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(342), ack => ptr_deref_1062_store_0_req_0); -- 
    maxPool4_cp_element_group_342: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_342"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(337) & maxPool4_CP_307_elements(341) & maxPool4_CP_307_elements(388) & maxPool4_CP_307_elements(344);
      gj_maxPool4_cp_element_group_342 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(342), clk => clk, reset => reset); --
    end block;
    -- CP-element group 343:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: marked-predecessors 
    -- CP-element group 343: 	345 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	345 
    -- CP-element group 343:  members (5) 
      -- CP-element group 343: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1062_Update/$entry
      -- CP-element group 343: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1062_Update/word_access_complete/$entry
      -- CP-element group 343: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1062_update_start_
      -- CP-element group 343: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1062_Update/word_access_complete/word_0/$entry
      -- CP-element group 343: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1062_Update/word_access_complete/word_0/cr
      -- 
    cr_1851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(343), ack => ptr_deref_1062_store_0_req_1); -- 
    maxPool4_cp_element_group_343: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_343"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_307_elements(345);
      gj_maxPool4_cp_element_group_343 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(343), clk => clk, reset => reset); --
    end block;
    -- CP-element group 344:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	342 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	389 
    -- CP-element group 344: marked-successors 
    -- CP-element group 344: 	335 
    -- CP-element group 344: 	339 
    -- CP-element group 344: 	342 
    -- CP-element group 344:  members (5) 
      -- CP-element group 344: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1062_sample_completed_
      -- CP-element group 344: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1062_Sample/$exit
      -- CP-element group 344: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1062_Sample/word_access_start/word_0/ra
      -- CP-element group 344: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1062_Sample/word_access_start/$exit
      -- CP-element group 344: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1062_Sample/word_access_start/word_0/$exit
      -- 
    ra_1841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 344_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1062_store_0_ack_0, ack => maxPool4_CP_307_elements(344)); -- 
    -- CP-element group 345:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	343 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	391 
    -- CP-element group 345: marked-successors 
    -- CP-element group 345: 	343 
    -- CP-element group 345:  members (5) 
      -- CP-element group 345: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1062_Update/$exit
      -- CP-element group 345: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1062_Update/word_access_complete/$exit
      -- CP-element group 345: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1062_update_completed_
      -- CP-element group 345: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1062_Update/word_access_complete/word_0/ca
      -- CP-element group 345: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1062_Update/word_access_complete/word_0/$exit
      -- 
    ca_1852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 345_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1062_store_0_ack_1, ack => maxPool4_CP_307_elements(345)); -- 
    -- CP-element group 346:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	350 
    -- CP-element group 346: marked-predecessors 
    -- CP-element group 346: 	351 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	351 
    -- CP-element group 346:  members (3) 
      -- CP-element group 346: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1082_request/$entry
      -- CP-element group 346: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1082_sample_start_
      -- CP-element group 346: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1082_request/req
      -- 
    req_1892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(346), ack => addr_of_1082_final_reg_req_0); -- 
    maxPool4_cp_element_group_346: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_346"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(350) & maxPool4_CP_307_elements(351);
      gj_maxPool4_cp_element_group_346 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(346), clk => clk, reset => reset); --
    end block;
    -- CP-element group 347:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	1 
    -- CP-element group 347: marked-predecessors 
    -- CP-element group 347: 	352 
    -- CP-element group 347: 	355 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	352 
    -- CP-element group 347:  members (3) 
      -- CP-element group 347: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1082_complete/$entry
      -- CP-element group 347: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1082_complete/req
      -- CP-element group 347: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1082_update_start_
      -- 
    req_1897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(347), ack => addr_of_1082_final_reg_req_1); -- 
    maxPool4_cp_element_group_347: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_347"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(1) & maxPool4_CP_307_elements(352) & maxPool4_CP_307_elements(355);
      gj_maxPool4_cp_element_group_347 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(347), clk => clk, reset => reset); --
    end block;
    -- CP-element group 348:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	1 
    -- CP-element group 348: marked-predecessors 
    -- CP-element group 348: 	350 
    -- CP-element group 348: 	351 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	350 
    -- CP-element group 348:  members (3) 
      -- CP-element group 348: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1081_final_index_sum_regn_update_start
      -- CP-element group 348: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1081_final_index_sum_regn_Update/req
      -- CP-element group 348: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1081_final_index_sum_regn_Update/$entry
      -- 
    req_1882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(348), ack => array_obj_ref_1081_index_offset_req_1); -- 
    maxPool4_cp_element_group_348: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_348"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(1) & maxPool4_CP_307_elements(350) & maxPool4_CP_307_elements(351);
      gj_maxPool4_cp_element_group_348 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(348), clk => clk, reset => reset); --
    end block;
    -- CP-element group 349:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	1 
    -- CP-element group 349: successors 
    -- CP-element group 349: 	391 
    -- CP-element group 349: marked-successors 
    -- CP-element group 349: 	2 
    -- CP-element group 349:  members (3) 
      -- CP-element group 349: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1081_final_index_sum_regn_Sample/$exit
      -- CP-element group 349: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1081_final_index_sum_regn_Sample/ack
      -- CP-element group 349: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1081_final_index_sum_regn_sample_complete
      -- 
    ack_1878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 349_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1081_index_offset_ack_0, ack => maxPool4_CP_307_elements(349)); -- 
    -- CP-element group 350:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	348 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	346 
    -- CP-element group 350: marked-successors 
    -- CP-element group 350: 	348 
    -- CP-element group 350:  members (8) 
      -- CP-element group 350: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1081_root_address_calculated
      -- CP-element group 350: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1081_final_index_sum_regn_Update/ack
      -- CP-element group 350: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1081_final_index_sum_regn_Update/$exit
      -- CP-element group 350: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1081_base_plus_offset/sum_rename_ack
      -- CP-element group 350: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1081_base_plus_offset/sum_rename_req
      -- CP-element group 350: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1081_base_plus_offset/$exit
      -- CP-element group 350: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1081_base_plus_offset/$entry
      -- CP-element group 350: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1081_offset_calculated
      -- 
    ack_1883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 350_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1081_index_offset_ack_1, ack => maxPool4_CP_307_elements(350)); -- 
    -- CP-element group 351:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	346 
    -- CP-element group 351: successors 
    -- CP-element group 351: marked-successors 
    -- CP-element group 351: 	346 
    -- CP-element group 351: 	348 
    -- CP-element group 351:  members (3) 
      -- CP-element group 351: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1082_request/ack
      -- CP-element group 351: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1082_request/$exit
      -- CP-element group 351: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1082_sample_completed_
      -- 
    ack_1893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 351_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1082_final_reg_ack_0, ack => maxPool4_CP_307_elements(351)); -- 
    -- CP-element group 352:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	347 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	353 
    -- CP-element group 352: marked-successors 
    -- CP-element group 352: 	347 
    -- CP-element group 352:  members (3) 
      -- CP-element group 352: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1082_complete/$exit
      -- CP-element group 352: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1082_complete/ack
      -- CP-element group 352: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1082_update_completed_
      -- 
    ack_1898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1082_final_reg_ack_1, ack => maxPool4_CP_307_elements(352)); -- 
    -- CP-element group 353:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	352 
    -- CP-element group 353: marked-predecessors 
    -- CP-element group 353: 	355 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	355 
    -- CP-element group 353:  members (3) 
      -- CP-element group 353: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1086_sample_start_
      -- CP-element group 353: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1086_Sample/$entry
      -- CP-element group 353: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1086_Sample/req
      -- 
    req_1906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(353), ack => W_myptr7_1078_delayed_8_0_1084_inst_req_0); -- 
    maxPool4_cp_element_group_353: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_353"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(352) & maxPool4_CP_307_elements(355);
      gj_maxPool4_cp_element_group_353 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(353), clk => clk, reset => reset); --
    end block;
    -- CP-element group 354:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: marked-predecessors 
    -- CP-element group 354: 	356 
    -- CP-element group 354: 	363 
    -- CP-element group 354: successors 
    -- CP-element group 354: 	356 
    -- CP-element group 354:  members (3) 
      -- CP-element group 354: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1086_update_start_
      -- CP-element group 354: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1086_Update/$entry
      -- CP-element group 354: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1086_Update/req
      -- 
    req_1911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(354), ack => W_myptr7_1078_delayed_8_0_1084_inst_req_1); -- 
    maxPool4_cp_element_group_354: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_354"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(356) & maxPool4_CP_307_elements(363);
      gj_maxPool4_cp_element_group_354 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(354), clk => clk, reset => reset); --
    end block;
    -- CP-element group 355:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	353 
    -- CP-element group 355: successors 
    -- CP-element group 355: marked-successors 
    -- CP-element group 355: 	347 
    -- CP-element group 355: 	353 
    -- CP-element group 355:  members (3) 
      -- CP-element group 355: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1086_sample_completed_
      -- CP-element group 355: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1086_Sample/$exit
      -- CP-element group 355: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1086_Sample/ack
      -- 
    ack_1907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 355_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_myptr7_1078_delayed_8_0_1084_inst_ack_0, ack => maxPool4_CP_307_elements(355)); -- 
    -- CP-element group 356:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	354 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	361 
    -- CP-element group 356: marked-successors 
    -- CP-element group 356: 	354 
    -- CP-element group 356:  members (19) 
      -- CP-element group 356: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1086_update_completed_
      -- CP-element group 356: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1086_Update/$exit
      -- CP-element group 356: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1086_Update/ack
      -- CP-element group 356: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1088_base_address_calculated
      -- CP-element group 356: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1088_word_address_calculated
      -- CP-element group 356: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1088_root_address_calculated
      -- CP-element group 356: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1088_base_address_resized
      -- CP-element group 356: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1088_base_addr_resize/$entry
      -- CP-element group 356: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1088_base_addr_resize/$exit
      -- CP-element group 356: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1088_base_addr_resize/base_resize_req
      -- CP-element group 356: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1088_base_addr_resize/base_resize_ack
      -- CP-element group 356: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1088_base_plus_offset/$entry
      -- CP-element group 356: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1088_base_plus_offset/$exit
      -- CP-element group 356: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1088_base_plus_offset/sum_rename_req
      -- CP-element group 356: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1088_base_plus_offset/sum_rename_ack
      -- CP-element group 356: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1088_word_addrgen/$entry
      -- CP-element group 356: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1088_word_addrgen/$exit
      -- CP-element group 356: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1088_word_addrgen/root_register_req
      -- CP-element group 356: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1088_word_addrgen/root_register_ack
      -- 
    ack_1912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 356_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_myptr7_1078_delayed_8_0_1084_inst_ack_1, ack => maxPool4_CP_307_elements(356)); -- 
    -- CP-element group 357:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	87 
    -- CP-element group 357: 	91 
    -- CP-element group 357: 	95 
    -- CP-element group 357: 	99 
    -- CP-element group 357: 	151 
    -- CP-element group 357: 	155 
    -- CP-element group 357: 	159 
    -- CP-element group 357: 	163 
    -- CP-element group 357: 	215 
    -- CP-element group 357: 	219 
    -- CP-element group 357: 	223 
    -- CP-element group 357: 	227 
    -- CP-element group 357: 	279 
    -- CP-element group 357: 	283 
    -- CP-element group 357: 	287 
    -- CP-element group 357: 	291 
    -- CP-element group 357: marked-predecessors 
    -- CP-element group 357: 	359 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	359 
    -- CP-element group 357:  members (3) 
      -- CP-element group 357: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1099_sample_start_
      -- CP-element group 357: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1099_Sample/$entry
      -- CP-element group 357: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1099_Sample/rr
      -- 
    rr_1920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(357), ack => CONCAT_u32_u64_1099_inst_req_0); -- 
    maxPool4_cp_element_group_357: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 1);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_357"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(87) & maxPool4_CP_307_elements(91) & maxPool4_CP_307_elements(95) & maxPool4_CP_307_elements(99) & maxPool4_CP_307_elements(151) & maxPool4_CP_307_elements(155) & maxPool4_CP_307_elements(159) & maxPool4_CP_307_elements(163) & maxPool4_CP_307_elements(215) & maxPool4_CP_307_elements(219) & maxPool4_CP_307_elements(223) & maxPool4_CP_307_elements(227) & maxPool4_CP_307_elements(279) & maxPool4_CP_307_elements(283) & maxPool4_CP_307_elements(287) & maxPool4_CP_307_elements(291) & maxPool4_CP_307_elements(359);
      gj_maxPool4_cp_element_group_357 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(357), clk => clk, reset => reset); --
    end block;
    -- CP-element group 358:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: marked-predecessors 
    -- CP-element group 358: 	360 
    -- CP-element group 358: 	363 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	360 
    -- CP-element group 358:  members (3) 
      -- CP-element group 358: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1099_update_start_
      -- CP-element group 358: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1099_Update/$entry
      -- CP-element group 358: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1099_Update/cr
      -- 
    cr_1925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(358), ack => CONCAT_u32_u64_1099_inst_req_1); -- 
    maxPool4_cp_element_group_358: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_358"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(360) & maxPool4_CP_307_elements(363);
      gj_maxPool4_cp_element_group_358 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(358), clk => clk, reset => reset); --
    end block;
    -- CP-element group 359:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	357 
    -- CP-element group 359: successors 
    -- CP-element group 359: marked-successors 
    -- CP-element group 359: 	85 
    -- CP-element group 359: 	89 
    -- CP-element group 359: 	93 
    -- CP-element group 359: 	97 
    -- CP-element group 359: 	149 
    -- CP-element group 359: 	153 
    -- CP-element group 359: 	157 
    -- CP-element group 359: 	161 
    -- CP-element group 359: 	213 
    -- CP-element group 359: 	217 
    -- CP-element group 359: 	221 
    -- CP-element group 359: 	225 
    -- CP-element group 359: 	277 
    -- CP-element group 359: 	281 
    -- CP-element group 359: 	285 
    -- CP-element group 359: 	289 
    -- CP-element group 359: 	357 
    -- CP-element group 359:  members (3) 
      -- CP-element group 359: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1099_sample_completed_
      -- CP-element group 359: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1099_Sample/$exit
      -- CP-element group 359: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1099_Sample/ra
      -- 
    ra_1921_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 359_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_1099_inst_ack_0, ack => maxPool4_CP_307_elements(359)); -- 
    -- CP-element group 360:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	358 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	361 
    -- CP-element group 360: marked-successors 
    -- CP-element group 360: 	358 
    -- CP-element group 360:  members (3) 
      -- CP-element group 360: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1099_update_completed_
      -- CP-element group 360: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1099_Update/$exit
      -- CP-element group 360: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1099_Update/ca
      -- 
    ca_1926_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 360_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_1099_inst_ack_1, ack => maxPool4_CP_307_elements(360)); -- 
    -- CP-element group 361:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	356 
    -- CP-element group 361: 	360 
    -- CP-element group 361: 	389 
    -- CP-element group 361: marked-predecessors 
    -- CP-element group 361: 	363 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	363 
    -- CP-element group 361:  members (9) 
      -- CP-element group 361: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1088_sample_start_
      -- CP-element group 361: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1088_Sample/$entry
      -- CP-element group 361: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1088_Sample/ptr_deref_1088_Split/$entry
      -- CP-element group 361: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1088_Sample/ptr_deref_1088_Split/$exit
      -- CP-element group 361: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1088_Sample/ptr_deref_1088_Split/split_req
      -- CP-element group 361: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1088_Sample/ptr_deref_1088_Split/split_ack
      -- CP-element group 361: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1088_Sample/word_access_start/$entry
      -- CP-element group 361: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1088_Sample/word_access_start/word_0/$entry
      -- CP-element group 361: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1088_Sample/word_access_start/word_0/rr
      -- 
    rr_1964_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1964_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(361), ack => ptr_deref_1088_store_0_req_0); -- 
    maxPool4_cp_element_group_361: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_361"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(356) & maxPool4_CP_307_elements(360) & maxPool4_CP_307_elements(389) & maxPool4_CP_307_elements(363);
      gj_maxPool4_cp_element_group_361 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(361), clk => clk, reset => reset); --
    end block;
    -- CP-element group 362:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: marked-predecessors 
    -- CP-element group 362: 	364 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	364 
    -- CP-element group 362:  members (5) 
      -- CP-element group 362: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1088_update_start_
      -- CP-element group 362: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1088_Update/$entry
      -- CP-element group 362: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1088_Update/word_access_complete/$entry
      -- CP-element group 362: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1088_Update/word_access_complete/word_0/$entry
      -- CP-element group 362: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1088_Update/word_access_complete/word_0/cr
      -- 
    cr_1975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(362), ack => ptr_deref_1088_store_0_req_1); -- 
    maxPool4_cp_element_group_362: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_362"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_307_elements(364);
      gj_maxPool4_cp_element_group_362 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(362), clk => clk, reset => reset); --
    end block;
    -- CP-element group 363:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	361 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	390 
    -- CP-element group 363: marked-successors 
    -- CP-element group 363: 	354 
    -- CP-element group 363: 	358 
    -- CP-element group 363: 	361 
    -- CP-element group 363:  members (5) 
      -- CP-element group 363: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1088_sample_completed_
      -- CP-element group 363: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1088_Sample/$exit
      -- CP-element group 363: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1088_Sample/word_access_start/$exit
      -- CP-element group 363: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1088_Sample/word_access_start/word_0/$exit
      -- CP-element group 363: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1088_Sample/word_access_start/word_0/ra
      -- 
    ra_1965_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 363_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1088_store_0_ack_0, ack => maxPool4_CP_307_elements(363)); -- 
    -- CP-element group 364:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	362 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	391 
    -- CP-element group 364: marked-successors 
    -- CP-element group 364: 	362 
    -- CP-element group 364:  members (5) 
      -- CP-element group 364: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1088_update_completed_
      -- CP-element group 364: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1088_Update/$exit
      -- CP-element group 364: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1088_Update/word_access_complete/$exit
      -- CP-element group 364: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1088_Update/word_access_complete/word_0/$exit
      -- CP-element group 364: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1088_Update/word_access_complete/word_0/ca
      -- 
    ca_1976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 364_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1088_store_0_ack_1, ack => maxPool4_CP_307_elements(364)); -- 
    -- CP-element group 365:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	369 
    -- CP-element group 365: marked-predecessors 
    -- CP-element group 365: 	370 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	370 
    -- CP-element group 365:  members (3) 
      -- CP-element group 365: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1108_sample_start_
      -- CP-element group 365: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1108_request/$entry
      -- CP-element group 365: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1108_request/req
      -- 
    req_2016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(365), ack => addr_of_1108_final_reg_req_0); -- 
    maxPool4_cp_element_group_365: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_365"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(369) & maxPool4_CP_307_elements(370);
      gj_maxPool4_cp_element_group_365 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(365), clk => clk, reset => reset); --
    end block;
    -- CP-element group 366:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	1 
    -- CP-element group 366: marked-predecessors 
    -- CP-element group 366: 	371 
    -- CP-element group 366: 	374 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	371 
    -- CP-element group 366:  members (3) 
      -- CP-element group 366: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1108_update_start_
      -- CP-element group 366: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1108_complete/$entry
      -- CP-element group 366: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1108_complete/req
      -- 
    req_2021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(366), ack => addr_of_1108_final_reg_req_1); -- 
    maxPool4_cp_element_group_366: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_366"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(1) & maxPool4_CP_307_elements(371) & maxPool4_CP_307_elements(374);
      gj_maxPool4_cp_element_group_366 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(366), clk => clk, reset => reset); --
    end block;
    -- CP-element group 367:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	1 
    -- CP-element group 367: marked-predecessors 
    -- CP-element group 367: 	369 
    -- CP-element group 367: 	370 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	369 
    -- CP-element group 367:  members (3) 
      -- CP-element group 367: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1107_final_index_sum_regn_update_start
      -- CP-element group 367: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1107_final_index_sum_regn_Update/$entry
      -- CP-element group 367: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1107_final_index_sum_regn_Update/req
      -- 
    req_2006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(367), ack => array_obj_ref_1107_index_offset_req_1); -- 
    maxPool4_cp_element_group_367: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_367"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(1) & maxPool4_CP_307_elements(369) & maxPool4_CP_307_elements(370);
      gj_maxPool4_cp_element_group_367 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(367), clk => clk, reset => reset); --
    end block;
    -- CP-element group 368:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	1 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	391 
    -- CP-element group 368: marked-successors 
    -- CP-element group 368: 	2 
    -- CP-element group 368:  members (3) 
      -- CP-element group 368: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1107_final_index_sum_regn_sample_complete
      -- CP-element group 368: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1107_final_index_sum_regn_Sample/$exit
      -- CP-element group 368: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1107_final_index_sum_regn_Sample/ack
      -- 
    ack_2002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 368_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1107_index_offset_ack_0, ack => maxPool4_CP_307_elements(368)); -- 
    -- CP-element group 369:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	367 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	365 
    -- CP-element group 369: marked-successors 
    -- CP-element group 369: 	367 
    -- CP-element group 369:  members (8) 
      -- CP-element group 369: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1107_root_address_calculated
      -- CP-element group 369: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1107_offset_calculated
      -- CP-element group 369: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1107_final_index_sum_regn_Update/$exit
      -- CP-element group 369: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1107_final_index_sum_regn_Update/ack
      -- CP-element group 369: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1107_base_plus_offset/$entry
      -- CP-element group 369: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1107_base_plus_offset/$exit
      -- CP-element group 369: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1107_base_plus_offset/sum_rename_req
      -- CP-element group 369: 	 assign_stmt_89_to_assign_stmt_1130/array_obj_ref_1107_base_plus_offset/sum_rename_ack
      -- 
    ack_2007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 369_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1107_index_offset_ack_1, ack => maxPool4_CP_307_elements(369)); -- 
    -- CP-element group 370:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	365 
    -- CP-element group 370: successors 
    -- CP-element group 370: marked-successors 
    -- CP-element group 370: 	365 
    -- CP-element group 370: 	367 
    -- CP-element group 370:  members (3) 
      -- CP-element group 370: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1108_sample_completed_
      -- CP-element group 370: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1108_request/$exit
      -- CP-element group 370: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1108_request/ack
      -- 
    ack_2017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 370_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1108_final_reg_ack_0, ack => maxPool4_CP_307_elements(370)); -- 
    -- CP-element group 371:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	366 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	372 
    -- CP-element group 371: marked-successors 
    -- CP-element group 371: 	366 
    -- CP-element group 371:  members (3) 
      -- CP-element group 371: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1108_update_completed_
      -- CP-element group 371: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1108_complete/$exit
      -- CP-element group 371: 	 assign_stmt_89_to_assign_stmt_1130/addr_of_1108_complete/ack
      -- 
    ack_2022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 371_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1108_final_reg_ack_1, ack => maxPool4_CP_307_elements(371)); -- 
    -- CP-element group 372:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	371 
    -- CP-element group 372: marked-predecessors 
    -- CP-element group 372: 	374 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	374 
    -- CP-element group 372:  members (3) 
      -- CP-element group 372: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1112_sample_start_
      -- CP-element group 372: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1112_Sample/$entry
      -- CP-element group 372: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1112_Sample/req
      -- 
    req_2030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(372), ack => W_myptr8_1101_delayed_8_0_1110_inst_req_0); -- 
    maxPool4_cp_element_group_372: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_372"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(371) & maxPool4_CP_307_elements(374);
      gj_maxPool4_cp_element_group_372 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(372), clk => clk, reset => reset); --
    end block;
    -- CP-element group 373:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: marked-predecessors 
    -- CP-element group 373: 	375 
    -- CP-element group 373: 	382 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	375 
    -- CP-element group 373:  members (3) 
      -- CP-element group 373: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1112_update_start_
      -- CP-element group 373: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1112_Update/$entry
      -- CP-element group 373: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1112_Update/req
      -- 
    req_2035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(373), ack => W_myptr8_1101_delayed_8_0_1110_inst_req_1); -- 
    maxPool4_cp_element_group_373: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_373"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(375) & maxPool4_CP_307_elements(382);
      gj_maxPool4_cp_element_group_373 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(373), clk => clk, reset => reset); --
    end block;
    -- CP-element group 374:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	372 
    -- CP-element group 374: successors 
    -- CP-element group 374: marked-successors 
    -- CP-element group 374: 	366 
    -- CP-element group 374: 	372 
    -- CP-element group 374:  members (3) 
      -- CP-element group 374: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1112_sample_completed_
      -- CP-element group 374: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1112_Sample/$exit
      -- CP-element group 374: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1112_Sample/ack
      -- 
    ack_2031_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 374_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_myptr8_1101_delayed_8_0_1110_inst_ack_0, ack => maxPool4_CP_307_elements(374)); -- 
    -- CP-element group 375:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	373 
    -- CP-element group 375: successors 
    -- CP-element group 375: 	380 
    -- CP-element group 375: marked-successors 
    -- CP-element group 375: 	373 
    -- CP-element group 375:  members (19) 
      -- CP-element group 375: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1112_update_completed_
      -- CP-element group 375: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1112_Update/$exit
      -- CP-element group 375: 	 assign_stmt_89_to_assign_stmt_1130/assign_stmt_1112_Update/ack
      -- CP-element group 375: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1114_base_address_calculated
      -- CP-element group 375: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1114_word_address_calculated
      -- CP-element group 375: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1114_root_address_calculated
      -- CP-element group 375: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1114_base_address_resized
      -- CP-element group 375: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1114_base_addr_resize/$entry
      -- CP-element group 375: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1114_base_addr_resize/$exit
      -- CP-element group 375: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1114_base_addr_resize/base_resize_req
      -- CP-element group 375: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1114_base_addr_resize/base_resize_ack
      -- CP-element group 375: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1114_base_plus_offset/$entry
      -- CP-element group 375: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1114_base_plus_offset/$exit
      -- CP-element group 375: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1114_base_plus_offset/sum_rename_req
      -- CP-element group 375: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1114_base_plus_offset/sum_rename_ack
      -- CP-element group 375: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1114_word_addrgen/$entry
      -- CP-element group 375: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1114_word_addrgen/$exit
      -- CP-element group 375: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1114_word_addrgen/root_register_req
      -- CP-element group 375: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1114_word_addrgen/root_register_ack
      -- 
    ack_2036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 375_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_myptr8_1101_delayed_8_0_1110_inst_ack_1, ack => maxPool4_CP_307_elements(375)); -- 
    -- CP-element group 376:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	103 
    -- CP-element group 376: 	107 
    -- CP-element group 376: 	111 
    -- CP-element group 376: 	115 
    -- CP-element group 376: 	167 
    -- CP-element group 376: 	171 
    -- CP-element group 376: 	175 
    -- CP-element group 376: 	179 
    -- CP-element group 376: 	231 
    -- CP-element group 376: 	235 
    -- CP-element group 376: 	239 
    -- CP-element group 376: 	243 
    -- CP-element group 376: 	295 
    -- CP-element group 376: 	299 
    -- CP-element group 376: 	303 
    -- CP-element group 376: 	307 
    -- CP-element group 376: marked-predecessors 
    -- CP-element group 376: 	378 
    -- CP-element group 376: successors 
    -- CP-element group 376: 	378 
    -- CP-element group 376:  members (3) 
      -- CP-element group 376: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1125_sample_start_
      -- CP-element group 376: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1125_Sample/$entry
      -- CP-element group 376: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1125_Sample/rr
      -- 
    rr_2044_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2044_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(376), ack => CONCAT_u32_u64_1125_inst_req_0); -- 
    maxPool4_cp_element_group_376: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 1);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_376"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(103) & maxPool4_CP_307_elements(107) & maxPool4_CP_307_elements(111) & maxPool4_CP_307_elements(115) & maxPool4_CP_307_elements(167) & maxPool4_CP_307_elements(171) & maxPool4_CP_307_elements(175) & maxPool4_CP_307_elements(179) & maxPool4_CP_307_elements(231) & maxPool4_CP_307_elements(235) & maxPool4_CP_307_elements(239) & maxPool4_CP_307_elements(243) & maxPool4_CP_307_elements(295) & maxPool4_CP_307_elements(299) & maxPool4_CP_307_elements(303) & maxPool4_CP_307_elements(307) & maxPool4_CP_307_elements(378);
      gj_maxPool4_cp_element_group_376 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(376), clk => clk, reset => reset); --
    end block;
    -- CP-element group 377:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: marked-predecessors 
    -- CP-element group 377: 	379 
    -- CP-element group 377: 	382 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	379 
    -- CP-element group 377:  members (3) 
      -- CP-element group 377: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1125_update_start_
      -- CP-element group 377: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1125_Update/$entry
      -- CP-element group 377: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1125_Update/cr
      -- 
    cr_2049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(377), ack => CONCAT_u32_u64_1125_inst_req_1); -- 
    maxPool4_cp_element_group_377: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_377"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(379) & maxPool4_CP_307_elements(382);
      gj_maxPool4_cp_element_group_377 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(377), clk => clk, reset => reset); --
    end block;
    -- CP-element group 378:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	376 
    -- CP-element group 378: successors 
    -- CP-element group 378: marked-successors 
    -- CP-element group 378: 	101 
    -- CP-element group 378: 	105 
    -- CP-element group 378: 	109 
    -- CP-element group 378: 	113 
    -- CP-element group 378: 	165 
    -- CP-element group 378: 	169 
    -- CP-element group 378: 	173 
    -- CP-element group 378: 	177 
    -- CP-element group 378: 	229 
    -- CP-element group 378: 	233 
    -- CP-element group 378: 	237 
    -- CP-element group 378: 	241 
    -- CP-element group 378: 	293 
    -- CP-element group 378: 	297 
    -- CP-element group 378: 	301 
    -- CP-element group 378: 	305 
    -- CP-element group 378: 	376 
    -- CP-element group 378:  members (3) 
      -- CP-element group 378: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1125_sample_completed_
      -- CP-element group 378: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1125_Sample/$exit
      -- CP-element group 378: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1125_Sample/ra
      -- 
    ra_2045_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 378_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_1125_inst_ack_0, ack => maxPool4_CP_307_elements(378)); -- 
    -- CP-element group 379:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	377 
    -- CP-element group 379: successors 
    -- CP-element group 379: 	380 
    -- CP-element group 379: marked-successors 
    -- CP-element group 379: 	377 
    -- CP-element group 379:  members (3) 
      -- CP-element group 379: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1125_update_completed_
      -- CP-element group 379: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1125_Update/$exit
      -- CP-element group 379: 	 assign_stmt_89_to_assign_stmt_1130/CONCAT_u32_u64_1125_Update/ca
      -- 
    ca_2050_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 379_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_1125_inst_ack_1, ack => maxPool4_CP_307_elements(379)); -- 
    -- CP-element group 380:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	375 
    -- CP-element group 380: 	379 
    -- CP-element group 380: 	390 
    -- CP-element group 380: marked-predecessors 
    -- CP-element group 380: 	382 
    -- CP-element group 380: successors 
    -- CP-element group 380: 	382 
    -- CP-element group 380:  members (9) 
      -- CP-element group 380: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1114_sample_start_
      -- CP-element group 380: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1114_Sample/$entry
      -- CP-element group 380: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1114_Sample/ptr_deref_1114_Split/$entry
      -- CP-element group 380: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1114_Sample/ptr_deref_1114_Split/$exit
      -- CP-element group 380: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1114_Sample/ptr_deref_1114_Split/split_req
      -- CP-element group 380: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1114_Sample/ptr_deref_1114_Split/split_ack
      -- CP-element group 380: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1114_Sample/word_access_start/$entry
      -- CP-element group 380: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1114_Sample/word_access_start/word_0/$entry
      -- CP-element group 380: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1114_Sample/word_access_start/word_0/rr
      -- 
    rr_2088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(380), ack => ptr_deref_1114_store_0_req_0); -- 
    maxPool4_cp_element_group_380: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_380"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(375) & maxPool4_CP_307_elements(379) & maxPool4_CP_307_elements(390) & maxPool4_CP_307_elements(382);
      gj_maxPool4_cp_element_group_380 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(380), clk => clk, reset => reset); --
    end block;
    -- CP-element group 381:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: marked-predecessors 
    -- CP-element group 381: 	383 
    -- CP-element group 381: successors 
    -- CP-element group 381: 	383 
    -- CP-element group 381:  members (5) 
      -- CP-element group 381: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1114_update_start_
      -- CP-element group 381: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1114_Update/$entry
      -- CP-element group 381: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1114_Update/word_access_complete/$entry
      -- CP-element group 381: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1114_Update/word_access_complete/word_0/$entry
      -- CP-element group 381: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1114_Update/word_access_complete/word_0/cr
      -- 
    cr_2099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(381), ack => ptr_deref_1114_store_0_req_1); -- 
    maxPool4_cp_element_group_381: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_381"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_307_elements(383);
      gj_maxPool4_cp_element_group_381 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(381), clk => clk, reset => reset); --
    end block;
    -- CP-element group 382:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	380 
    -- CP-element group 382: successors 
    -- CP-element group 382: 	391 
    -- CP-element group 382: marked-successors 
    -- CP-element group 382: 	323 
    -- CP-element group 382: 	373 
    -- CP-element group 382: 	377 
    -- CP-element group 382: 	380 
    -- CP-element group 382:  members (6) 
      -- CP-element group 382: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1114_sample_completed_
      -- CP-element group 382: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1114_Sample/$exit
      -- CP-element group 382: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1114_Sample/word_access_start/$exit
      -- CP-element group 382: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1114_Sample/word_access_start/word_0/$exit
      -- CP-element group 382: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1114_Sample/word_access_start/word_0/ra
      -- CP-element group 382: 	 assign_stmt_89_to_assign_stmt_1130/ring_reenable_memory_space_0
      -- 
    ra_2089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 382_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1114_store_0_ack_0, ack => maxPool4_CP_307_elements(382)); -- 
    -- CP-element group 383:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	381 
    -- CP-element group 383: successors 
    -- CP-element group 383: 	391 
    -- CP-element group 383: marked-successors 
    -- CP-element group 383: 	381 
    -- CP-element group 383:  members (5) 
      -- CP-element group 383: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1114_update_completed_
      -- CP-element group 383: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1114_Update/$exit
      -- CP-element group 383: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1114_Update/word_access_complete/$exit
      -- CP-element group 383: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1114_Update/word_access_complete/word_0/$exit
      -- CP-element group 383: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1114_Update/word_access_complete/word_0/ca
      -- 
    ca_2100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 383_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1114_store_0_ack_1, ack => maxPool4_CP_307_elements(383)); -- 
    -- CP-element group 384:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	55 
    -- CP-element group 384: 	119 
    -- CP-element group 384: 	183 
    -- CP-element group 384: 	247 
    -- CP-element group 384: marked-predecessors 
    -- CP-element group 384: 	386 
    -- CP-element group 384: successors 
    -- CP-element group 384: 	386 
    -- CP-element group 384:  members (3) 
      -- CP-element group 384: 	 assign_stmt_89_to_assign_stmt_1130/type_cast_1129_sample_start_
      -- CP-element group 384: 	 assign_stmt_89_to_assign_stmt_1130/type_cast_1129_Sample/$entry
      -- CP-element group 384: 	 assign_stmt_89_to_assign_stmt_1130/type_cast_1129_Sample/rr
      -- 
    rr_2108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(384), ack => type_cast_1129_inst_req_0); -- 
    maxPool4_cp_element_group_384: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_384"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(55) & maxPool4_CP_307_elements(119) & maxPool4_CP_307_elements(183) & maxPool4_CP_307_elements(247) & maxPool4_CP_307_elements(386);
      gj_maxPool4_cp_element_group_384 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(384), clk => clk, reset => reset); --
    end block;
    -- CP-element group 385:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	7 
    -- CP-element group 385: marked-predecessors 
    -- CP-element group 385: 	387 
    -- CP-element group 385: successors 
    -- CP-element group 385: 	387 
    -- CP-element group 385:  members (3) 
      -- CP-element group 385: 	 assign_stmt_89_to_assign_stmt_1130/type_cast_1129_update_start_
      -- CP-element group 385: 	 assign_stmt_89_to_assign_stmt_1130/type_cast_1129_Update/$entry
      -- CP-element group 385: 	 assign_stmt_89_to_assign_stmt_1130/type_cast_1129_Update/cr
      -- 
    cr_2113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_307_elements(385), ack => type_cast_1129_inst_req_1); -- 
    maxPool4_cp_element_group_385: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_385"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(7) & maxPool4_CP_307_elements(387);
      gj_maxPool4_cp_element_group_385 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(385), clk => clk, reset => reset); --
    end block;
    -- CP-element group 386:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	384 
    -- CP-element group 386: successors 
    -- CP-element group 386: marked-successors 
    -- CP-element group 386: 	53 
    -- CP-element group 386: 	117 
    -- CP-element group 386: 	181 
    -- CP-element group 386: 	245 
    -- CP-element group 386: 	384 
    -- CP-element group 386:  members (3) 
      -- CP-element group 386: 	 assign_stmt_89_to_assign_stmt_1130/type_cast_1129_sample_completed_
      -- CP-element group 386: 	 assign_stmt_89_to_assign_stmt_1130/type_cast_1129_Sample/$exit
      -- CP-element group 386: 	 assign_stmt_89_to_assign_stmt_1130/type_cast_1129_Sample/ra
      -- 
    ra_2109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 386_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1129_inst_ack_0, ack => maxPool4_CP_307_elements(386)); -- 
    -- CP-element group 387:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	385 
    -- CP-element group 387: successors 
    -- CP-element group 387: 	391 
    -- CP-element group 387: marked-successors 
    -- CP-element group 387: 	385 
    -- CP-element group 387:  members (3) 
      -- CP-element group 387: 	 assign_stmt_89_to_assign_stmt_1130/type_cast_1129_update_completed_
      -- CP-element group 387: 	 assign_stmt_89_to_assign_stmt_1130/type_cast_1129_Update/$exit
      -- CP-element group 387: 	 assign_stmt_89_to_assign_stmt_1130/type_cast_1129_Update/ca
      -- 
    ca_2114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 387_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1129_inst_ack_1, ack => maxPool4_CP_307_elements(387)); -- 
    -- CP-element group 388:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: 	325 
    -- CP-element group 388: successors 
    -- CP-element group 388: 	342 
    -- CP-element group 388:  members (1) 
      -- CP-element group 388: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1036_ptr_deref_1062_delay
      -- 
    -- Element group maxPool4_CP_307_elements(388) is a control-delay.
    cp_element_388_delay: control_delay_element  generic map(name => " 388_delay", delay_value => 1)  port map(req => maxPool4_CP_307_elements(325), ack => maxPool4_CP_307_elements(388), clk => clk, reset =>reset);
    -- CP-element group 389:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	344 
    -- CP-element group 389: successors 
    -- CP-element group 389: 	361 
    -- CP-element group 389:  members (1) 
      -- CP-element group 389: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1062_ptr_deref_1088_delay
      -- 
    -- Element group maxPool4_CP_307_elements(389) is a control-delay.
    cp_element_389_delay: control_delay_element  generic map(name => " 389_delay", delay_value => 1)  port map(req => maxPool4_CP_307_elements(344), ack => maxPool4_CP_307_elements(389), clk => clk, reset =>reset);
    -- CP-element group 390:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: 	363 
    -- CP-element group 390: successors 
    -- CP-element group 390: 	380 
    -- CP-element group 390:  members (1) 
      -- CP-element group 390: 	 assign_stmt_89_to_assign_stmt_1130/ptr_deref_1088_ptr_deref_1114_delay
      -- 
    -- Element group maxPool4_CP_307_elements(390) is a control-delay.
    cp_element_390_delay: control_delay_element  generic map(name => " 390_delay", delay_value => 1)  port map(req => maxPool4_CP_307_elements(363), ack => maxPool4_CP_307_elements(390), clk => clk, reset =>reset);
    -- CP-element group 391:  join  transition  bypass  pipeline-parent 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: 	11 
    -- CP-element group 391: 	18 
    -- CP-element group 391: 	25 
    -- CP-element group 391: 	32 
    -- CP-element group 391: 	311 
    -- CP-element group 391: 	326 
    -- CP-element group 391: 	330 
    -- CP-element group 391: 	345 
    -- CP-element group 391: 	349 
    -- CP-element group 391: 	364 
    -- CP-element group 391: 	368 
    -- CP-element group 391: 	382 
    -- CP-element group 391: 	383 
    -- CP-element group 391: 	387 
    -- CP-element group 391: successors 
    -- CP-element group 391: 	398 
    -- CP-element group 391:  members (1) 
      -- CP-element group 391: 	 assign_stmt_89_to_assign_stmt_1130/$exit
      -- 
    maxPool4_cp_element_group_391: block -- 
      constant place_capacities: IntegerArray(0 to 13) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 15,11 => 15,12 => 15,13 => 15);
      constant place_markings: IntegerArray(0 to 13)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0);
      constant place_delays: IntegerArray(0 to 13) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_391"; 
      signal preds: BooleanArray(1 to 14); -- 
    begin -- 
      preds <= maxPool4_CP_307_elements(11) & maxPool4_CP_307_elements(18) & maxPool4_CP_307_elements(25) & maxPool4_CP_307_elements(32) & maxPool4_CP_307_elements(311) & maxPool4_CP_307_elements(326) & maxPool4_CP_307_elements(330) & maxPool4_CP_307_elements(345) & maxPool4_CP_307_elements(349) & maxPool4_CP_307_elements(364) & maxPool4_CP_307_elements(368) & maxPool4_CP_307_elements(382) & maxPool4_CP_307_elements(383) & maxPool4_CP_307_elements(387);
      gj_maxPool4_cp_element_group_391 : generic_join generic map(name => joinName, number_of_predecessors => 14, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_307_elements(391), clk => clk, reset => reset); --
    end block;
    -- CP-element group 392:  place  bypass  pipeline-parent 
    -- CP-element group 392: predecessors 
    -- CP-element group 392: 	2 
    -- CP-element group 392: successors 
    -- CP-element group 392:  members (1) 
      -- CP-element group 392: 	 addr_update_enable
      -- 
    maxPool4_CP_307_elements(392) <= maxPool4_CP_307_elements(2);
    -- CP-element group 393:  place  bypass  pipeline-parent 
    -- CP-element group 393: predecessors 
    -- CP-element group 393: 	3 
    -- CP-element group 393: successors 
    -- CP-element group 393:  members (1) 
      -- CP-element group 393: 	 addr1_update_enable
      -- 
    maxPool4_CP_307_elements(393) <= maxPool4_CP_307_elements(3);
    -- CP-element group 394:  place  bypass  pipeline-parent 
    -- CP-element group 394: predecessors 
    -- CP-element group 394: 	4 
    -- CP-element group 394: successors 
    -- CP-element group 394:  members (1) 
      -- CP-element group 394: 	 addr2_update_enable
      -- 
    maxPool4_CP_307_elements(394) <= maxPool4_CP_307_elements(4);
    -- CP-element group 395:  place  bypass  pipeline-parent 
    -- CP-element group 395: predecessors 
    -- CP-element group 395: 	5 
    -- CP-element group 395: successors 
    -- CP-element group 395:  members (1) 
      -- CP-element group 395: 	 addr3_update_enable
      -- 
    maxPool4_CP_307_elements(395) <= maxPool4_CP_307_elements(5);
    -- CP-element group 396:  place  bypass  pipeline-parent 
    -- CP-element group 396: predecessors 
    -- CP-element group 396: 	6 
    -- CP-element group 396: successors 
    -- CP-element group 396:  members (1) 
      -- CP-element group 396: 	 addr4_update_enable
      -- 
    maxPool4_CP_307_elements(396) <= maxPool4_CP_307_elements(6);
    -- CP-element group 397:  place  bypass  pipeline-parent 
    -- CP-element group 397: predecessors 
    -- CP-element group 397: successors 
    -- CP-element group 397: 	7 
    -- CP-element group 397:  members (1) 
      -- CP-element group 397: 	 output_update_enable
      -- 
    -- CP-element group 398:  transition  bypass  pipeline-parent 
    -- CP-element group 398: predecessors 
    -- CP-element group 398: 	391 
    -- CP-element group 398: successors 
    -- CP-element group 398:  members (1) 
      -- CP-element group 398: 	 $exit
      -- 
    maxPool4_CP_307_elements(398) <= maxPool4_CP_307_elements(391);
    --  hookup: inputs to control-path 
    maxPool4_CP_307_elements(397) <= output_update_enable;
    -- hookup: output from control-path 
    addr_update_enable <= maxPool4_CP_307_elements(392);
    addr1_update_enable <= maxPool4_CP_307_elements(393);
    addr2_update_enable <= maxPool4_CP_307_elements(394);
    addr3_update_enable <= maxPool4_CP_307_elements(395);
    addr4_update_enable <= maxPool4_CP_307_elements(396);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u32_u32_1054_resized : std_logic_vector(13 downto 0);
    signal ADD_u32_u32_1054_scaled : std_logic_vector(13 downto 0);
    signal ADD_u32_u32_1054_wire : std_logic_vector(31 downto 0);
    signal ADD_u32_u32_1080_resized : std_logic_vector(13 downto 0);
    signal ADD_u32_u32_1080_scaled : std_logic_vector(13 downto 0);
    signal ADD_u32_u32_1080_wire : std_logic_vector(31 downto 0);
    signal ADD_u32_u32_1106_resized : std_logic_vector(13 downto 0);
    signal ADD_u32_u32_1106_scaled : std_logic_vector(13 downto 0);
    signal ADD_u32_u32_1106_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_1041_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_1046_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_1067_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_1072_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_1093_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_1098_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_1119_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_1124_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u32_u64_1047_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u32_u64_1073_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u32_u64_1099_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u32_u64_1125_wire : std_logic_vector(63 downto 0);
    signal R_addr1_86_resized : std_logic_vector(13 downto 0);
    signal R_addr1_86_scaled : std_logic_vector(13 downto 0);
    signal R_addr2_93_resized : std_logic_vector(13 downto 0);
    signal R_addr2_93_scaled : std_logic_vector(13 downto 0);
    signal R_addr3_100_resized : std_logic_vector(13 downto 0);
    signal R_addr3_100_scaled : std_logic_vector(13 downto 0);
    signal R_addr4_107_resized : std_logic_vector(13 downto 0);
    signal R_addr4_107_scaled : std_logic_vector(13 downto 0);
    signal R_addr_1028_resized : std_logic_vector(13 downto 0);
    signal R_addr_1028_scaled : std_logic_vector(13 downto 0);
    signal SGT_i16_u1_1004_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1012_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1020_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_644_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_652_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_660_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_668_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_676_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_684_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_692_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_700_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_708_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_716_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_724_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_732_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_740_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_748_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_756_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_764_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_772_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_780_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_788_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_796_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_804_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_812_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_820_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_828_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_836_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_844_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_852_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_860_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_868_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_876_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_884_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_892_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_900_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_908_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_916_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_924_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_932_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_940_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_948_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_956_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_964_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_972_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_980_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_988_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_996_wire : std_logic_vector(0 downto 0);
    signal a110_424 : std_logic_vector(15 downto 0);
    signal a111_428 : std_logic_vector(15 downto 0);
    signal a112_432 : std_logic_vector(15 downto 0);
    signal a113_436 : std_logic_vector(15 downto 0);
    signal a114_440 : std_logic_vector(15 downto 0);
    signal a115_444 : std_logic_vector(15 downto 0);
    signal a116_448 : std_logic_vector(15 downto 0);
    signal a11_388 : std_logic_vector(15 downto 0);
    signal a12_392 : std_logic_vector(15 downto 0);
    signal a13_396 : std_logic_vector(15 downto 0);
    signal a14_400 : std_logic_vector(15 downto 0);
    signal a15_404 : std_logic_vector(15 downto 0);
    signal a16_408 : std_logic_vector(15 downto 0);
    signal a17_412 : std_logic_vector(15 downto 0);
    signal a18_416 : std_logic_vector(15 downto 0);
    signal a19_420 : std_logic_vector(15 downto 0);
    signal a210_488 : std_logic_vector(15 downto 0);
    signal a211_492 : std_logic_vector(15 downto 0);
    signal a212_496 : std_logic_vector(15 downto 0);
    signal a213_500 : std_logic_vector(15 downto 0);
    signal a214_504 : std_logic_vector(15 downto 0);
    signal a215_508 : std_logic_vector(15 downto 0);
    signal a216_512 : std_logic_vector(15 downto 0);
    signal a21_452 : std_logic_vector(15 downto 0);
    signal a22_456 : std_logic_vector(15 downto 0);
    signal a23_460 : std_logic_vector(15 downto 0);
    signal a24_464 : std_logic_vector(15 downto 0);
    signal a25_468 : std_logic_vector(15 downto 0);
    signal a26_472 : std_logic_vector(15 downto 0);
    signal a27_476 : std_logic_vector(15 downto 0);
    signal a28_480 : std_logic_vector(15 downto 0);
    signal a29_484 : std_logic_vector(15 downto 0);
    signal a310_552 : std_logic_vector(15 downto 0);
    signal a311_556 : std_logic_vector(15 downto 0);
    signal a312_560 : std_logic_vector(15 downto 0);
    signal a313_564 : std_logic_vector(15 downto 0);
    signal a314_568 : std_logic_vector(15 downto 0);
    signal a315_572 : std_logic_vector(15 downto 0);
    signal a316_576 : std_logic_vector(15 downto 0);
    signal a31_516 : std_logic_vector(15 downto 0);
    signal a32_520 : std_logic_vector(15 downto 0);
    signal a33_524 : std_logic_vector(15 downto 0);
    signal a34_528 : std_logic_vector(15 downto 0);
    signal a35_532 : std_logic_vector(15 downto 0);
    signal a36_536 : std_logic_vector(15 downto 0);
    signal a37_540 : std_logic_vector(15 downto 0);
    signal a38_544 : std_logic_vector(15 downto 0);
    signal a39_548 : std_logic_vector(15 downto 0);
    signal a410_616 : std_logic_vector(15 downto 0);
    signal a411_620 : std_logic_vector(15 downto 0);
    signal a412_624 : std_logic_vector(15 downto 0);
    signal a413_628 : std_logic_vector(15 downto 0);
    signal a414_632 : std_logic_vector(15 downto 0);
    signal a415_636 : std_logic_vector(15 downto 0);
    signal a416_640 : std_logic_vector(15 downto 0);
    signal a41_580 : std_logic_vector(15 downto 0);
    signal a42_584 : std_logic_vector(15 downto 0);
    signal a43_588 : std_logic_vector(15 downto 0);
    signal a44_592 : std_logic_vector(15 downto 0);
    signal a45_596 : std_logic_vector(15 downto 0);
    signal a46_600 : std_logic_vector(15 downto 0);
    signal a47_604 : std_logic_vector(15 downto 0);
    signal a48_608 : std_logic_vector(15 downto 0);
    signal a49_612 : std_logic_vector(15 downto 0);
    signal array_obj_ref_101_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_101_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_101_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_101_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_101_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_101_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1029_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1029_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1029_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1029_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1029_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1029_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1055_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1055_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1055_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1055_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1055_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1055_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1081_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1081_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1081_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1081_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1081_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1081_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_108_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_108_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_108_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_108_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_108_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_108_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1107_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1107_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1107_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1107_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1107_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1107_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_87_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_87_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_87_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_87_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_87_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_87_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_94_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_94_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_94_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_94_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_94_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_94_root_address : std_logic_vector(13 downto 0);
    signal c1_114 : std_logic_vector(255 downto 0);
    signal c2_118 : std_logic_vector(255 downto 0);
    signal c3_122 : std_logic_vector(255 downto 0);
    signal c4_126 : std_logic_vector(255 downto 0);
    signal konst_1053_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1079_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1105_wire_constant : std_logic_vector(31 downto 0);
    signal myptr1_89 : std_logic_vector(31 downto 0);
    signal myptr2_96 : std_logic_vector(31 downto 0);
    signal myptr3_103 : std_logic_vector(31 downto 0);
    signal myptr4_110 : std_logic_vector(31 downto 0);
    signal myptr5_1031 : std_logic_vector(31 downto 0);
    signal myptr5_1032_delayed_8_0_1034 : std_logic_vector(31 downto 0);
    signal myptr6_1055_delayed_8_0_1060 : std_logic_vector(31 downto 0);
    signal myptr6_1057 : std_logic_vector(31 downto 0);
    signal myptr7_1078_delayed_8_0_1086 : std_logic_vector(31 downto 0);
    signal myptr7_1083 : std_logic_vector(31 downto 0);
    signal myptr8_1101_delayed_8_0_1112 : std_logic_vector(31 downto 0);
    signal myptr8_1109 : std_logic_vector(31 downto 0);
    signal out10_880 : std_logic_vector(15 downto 0);
    signal out11_904 : std_logic_vector(15 downto 0);
    signal out12_928 : std_logic_vector(15 downto 0);
    signal out13_952 : std_logic_vector(15 downto 0);
    signal out14_976 : std_logic_vector(15 downto 0);
    signal out15_1000 : std_logic_vector(15 downto 0);
    signal out16_1024 : std_logic_vector(15 downto 0);
    signal out1_664 : std_logic_vector(15 downto 0);
    signal out2_688 : std_logic_vector(15 downto 0);
    signal out3_712 : std_logic_vector(15 downto 0);
    signal out4_736 : std_logic_vector(15 downto 0);
    signal out5_760 : std_logic_vector(15 downto 0);
    signal out6_784 : std_logic_vector(15 downto 0);
    signal out7_808 : std_logic_vector(15 downto 0);
    signal out8_832 : std_logic_vector(15 downto 0);
    signal out9_856 : std_logic_vector(15 downto 0);
    signal ptr_deref_1036_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1036_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1036_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1036_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1036_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1036_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1062_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1062_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1062_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1062_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1062_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1062_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1088_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1088_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1088_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1088_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1088_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1088_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1114_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1114_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1114_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1114_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1114_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1114_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_113_data_0 : std_logic_vector(255 downto 0);
    signal ptr_deref_113_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_113_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_113_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_113_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_117_data_0 : std_logic_vector(255 downto 0);
    signal ptr_deref_117_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_117_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_117_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_117_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_121_data_0 : std_logic_vector(255 downto 0);
    signal ptr_deref_121_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_121_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_121_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_121_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_125_data_0 : std_logic_vector(255 downto 0);
    signal ptr_deref_125_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_125_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_125_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_125_word_offset_0 : std_logic_vector(13 downto 0);
    signal sliced_v110_167 : std_logic_vector(15 downto 0);
    signal sliced_v111_171 : std_logic_vector(15 downto 0);
    signal sliced_v112_175 : std_logic_vector(15 downto 0);
    signal sliced_v113_179 : std_logic_vector(15 downto 0);
    signal sliced_v114_183 : std_logic_vector(15 downto 0);
    signal sliced_v115_187 : std_logic_vector(15 downto 0);
    signal sliced_v116_191 : std_logic_vector(15 downto 0);
    signal sliced_v11_131 : std_logic_vector(15 downto 0);
    signal sliced_v12_135 : std_logic_vector(15 downto 0);
    signal sliced_v13_139 : std_logic_vector(15 downto 0);
    signal sliced_v14_143 : std_logic_vector(15 downto 0);
    signal sliced_v15_147 : std_logic_vector(15 downto 0);
    signal sliced_v16_151 : std_logic_vector(15 downto 0);
    signal sliced_v17_155 : std_logic_vector(15 downto 0);
    signal sliced_v18_159 : std_logic_vector(15 downto 0);
    signal sliced_v19_163 : std_logic_vector(15 downto 0);
    signal sliced_v210_231 : std_logic_vector(15 downto 0);
    signal sliced_v211_235 : std_logic_vector(15 downto 0);
    signal sliced_v212_239 : std_logic_vector(15 downto 0);
    signal sliced_v213_243 : std_logic_vector(15 downto 0);
    signal sliced_v214_247 : std_logic_vector(15 downto 0);
    signal sliced_v215_251 : std_logic_vector(15 downto 0);
    signal sliced_v216_255 : std_logic_vector(15 downto 0);
    signal sliced_v21_195 : std_logic_vector(15 downto 0);
    signal sliced_v22_199 : std_logic_vector(15 downto 0);
    signal sliced_v23_203 : std_logic_vector(15 downto 0);
    signal sliced_v24_207 : std_logic_vector(15 downto 0);
    signal sliced_v25_211 : std_logic_vector(15 downto 0);
    signal sliced_v26_215 : std_logic_vector(15 downto 0);
    signal sliced_v27_219 : std_logic_vector(15 downto 0);
    signal sliced_v28_223 : std_logic_vector(15 downto 0);
    signal sliced_v29_227 : std_logic_vector(15 downto 0);
    signal sliced_v310_295 : std_logic_vector(15 downto 0);
    signal sliced_v311_299 : std_logic_vector(15 downto 0);
    signal sliced_v312_303 : std_logic_vector(15 downto 0);
    signal sliced_v313_307 : std_logic_vector(15 downto 0);
    signal sliced_v314_311 : std_logic_vector(15 downto 0);
    signal sliced_v315_315 : std_logic_vector(15 downto 0);
    signal sliced_v316_319 : std_logic_vector(15 downto 0);
    signal sliced_v31_259 : std_logic_vector(15 downto 0);
    signal sliced_v32_263 : std_logic_vector(15 downto 0);
    signal sliced_v33_267 : std_logic_vector(15 downto 0);
    signal sliced_v34_271 : std_logic_vector(15 downto 0);
    signal sliced_v35_275 : std_logic_vector(15 downto 0);
    signal sliced_v36_279 : std_logic_vector(15 downto 0);
    signal sliced_v37_283 : std_logic_vector(15 downto 0);
    signal sliced_v38_287 : std_logic_vector(15 downto 0);
    signal sliced_v39_291 : std_logic_vector(15 downto 0);
    signal sliced_v410_359 : std_logic_vector(15 downto 0);
    signal sliced_v411_363 : std_logic_vector(15 downto 0);
    signal sliced_v412_367 : std_logic_vector(15 downto 0);
    signal sliced_v413_371 : std_logic_vector(15 downto 0);
    signal sliced_v414_375 : std_logic_vector(15 downto 0);
    signal sliced_v415_379 : std_logic_vector(15 downto 0);
    signal sliced_v416_383 : std_logic_vector(15 downto 0);
    signal sliced_v41_323 : std_logic_vector(15 downto 0);
    signal sliced_v42_327 : std_logic_vector(15 downto 0);
    signal sliced_v43_331 : std_logic_vector(15 downto 0);
    signal sliced_v44_335 : std_logic_vector(15 downto 0);
    signal sliced_v45_339 : std_logic_vector(15 downto 0);
    signal sliced_v46_343 : std_logic_vector(15 downto 0);
    signal sliced_v47_347 : std_logic_vector(15 downto 0);
    signal sliced_v48_351 : std_logic_vector(15 downto 0);
    signal sliced_v49_355 : std_logic_vector(15 downto 0);
    signal t101_864 : std_logic_vector(15 downto 0);
    signal t102_872 : std_logic_vector(15 downto 0);
    signal t111_888 : std_logic_vector(15 downto 0);
    signal t112_896 : std_logic_vector(15 downto 0);
    signal t11_648 : std_logic_vector(15 downto 0);
    signal t121_912 : std_logic_vector(15 downto 0);
    signal t122_920 : std_logic_vector(15 downto 0);
    signal t12_656 : std_logic_vector(15 downto 0);
    signal t131_936 : std_logic_vector(15 downto 0);
    signal t132_944 : std_logic_vector(15 downto 0);
    signal t141_960 : std_logic_vector(15 downto 0);
    signal t142_968 : std_logic_vector(15 downto 0);
    signal t151_984 : std_logic_vector(15 downto 0);
    signal t152_992 : std_logic_vector(15 downto 0);
    signal t161_1008 : std_logic_vector(15 downto 0);
    signal t162_1016 : std_logic_vector(15 downto 0);
    signal t21_672 : std_logic_vector(15 downto 0);
    signal t22_680 : std_logic_vector(15 downto 0);
    signal t31_696 : std_logic_vector(15 downto 0);
    signal t32_704 : std_logic_vector(15 downto 0);
    signal t41_720 : std_logic_vector(15 downto 0);
    signal t42_728 : std_logic_vector(15 downto 0);
    signal t51_744 : std_logic_vector(15 downto 0);
    signal t52_752 : std_logic_vector(15 downto 0);
    signal t61_768 : std_logic_vector(15 downto 0);
    signal t62_776 : std_logic_vector(15 downto 0);
    signal t71_792 : std_logic_vector(15 downto 0);
    signal t72_800 : std_logic_vector(15 downto 0);
    signal t81_816 : std_logic_vector(15 downto 0);
    signal t82_824 : std_logic_vector(15 downto 0);
    signal t91_840 : std_logic_vector(15 downto 0);
    signal t92_848 : std_logic_vector(15 downto 0);
    signal type_cast_1038_wire : std_logic_vector(15 downto 0);
    signal type_cast_1040_wire : std_logic_vector(15 downto 0);
    signal type_cast_1043_wire : std_logic_vector(15 downto 0);
    signal type_cast_1045_wire : std_logic_vector(15 downto 0);
    signal type_cast_1064_wire : std_logic_vector(15 downto 0);
    signal type_cast_1066_wire : std_logic_vector(15 downto 0);
    signal type_cast_1069_wire : std_logic_vector(15 downto 0);
    signal type_cast_1071_wire : std_logic_vector(15 downto 0);
    signal type_cast_1090_wire : std_logic_vector(15 downto 0);
    signal type_cast_1092_wire : std_logic_vector(15 downto 0);
    signal type_cast_1095_wire : std_logic_vector(15 downto 0);
    signal type_cast_1097_wire : std_logic_vector(15 downto 0);
    signal type_cast_1116_wire : std_logic_vector(15 downto 0);
    signal type_cast_1118_wire : std_logic_vector(15 downto 0);
    signal type_cast_1121_wire : std_logic_vector(15 downto 0);
    signal type_cast_1123_wire : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_101_constant_part_of_offset <= "00000000000000";
    array_obj_ref_101_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_101_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_101_resized_base_address <= "00000000000000";
    array_obj_ref_1029_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1029_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1029_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1029_resized_base_address <= "00000000000000";
    array_obj_ref_1055_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1055_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1055_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1055_resized_base_address <= "00000000000000";
    array_obj_ref_1081_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1081_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1081_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1081_resized_base_address <= "00000000000000";
    array_obj_ref_108_constant_part_of_offset <= "00000000000000";
    array_obj_ref_108_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_108_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_108_resized_base_address <= "00000000000000";
    array_obj_ref_1107_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1107_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1107_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1107_resized_base_address <= "00000000000000";
    array_obj_ref_87_constant_part_of_offset <= "00000000000000";
    array_obj_ref_87_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_87_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_87_resized_base_address <= "00000000000000";
    array_obj_ref_94_constant_part_of_offset <= "00000000000000";
    array_obj_ref_94_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_94_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_94_resized_base_address <= "00000000000000";
    konst_1053_wire_constant <= "00000000000000000000000000000001";
    konst_1079_wire_constant <= "00000000000000000000000000000010";
    konst_1105_wire_constant <= "00000000000000000000000000000011";
    ptr_deref_1036_word_offset_0 <= "00000000000000";
    ptr_deref_1062_word_offset_0 <= "00000000000000";
    ptr_deref_1088_word_offset_0 <= "00000000000000";
    ptr_deref_1114_word_offset_0 <= "00000000000000";
    ptr_deref_113_word_offset_0 <= "00000000000000";
    ptr_deref_117_word_offset_0 <= "00000000000000";
    ptr_deref_121_word_offset_0 <= "00000000000000";
    ptr_deref_125_word_offset_0 <= "00000000000000";
    -- flow-through select operator MUX_1007_inst
    t161_1008 <= a116_448 when (SGT_i16_u1_1004_wire(0) /=  '0') else a216_512;
    -- flow-through select operator MUX_1015_inst
    t162_1016 <= a316_576 when (SGT_i16_u1_1012_wire(0) /=  '0') else a416_640;
    -- flow-through select operator MUX_1023_inst
    out16_1024 <= t161_1008 when (SGT_i16_u1_1020_wire(0) /=  '0') else t162_1016;
    -- flow-through select operator MUX_647_inst
    t11_648 <= a11_388 when (SGT_i16_u1_644_wire(0) /=  '0') else a21_452;
    -- flow-through select operator MUX_655_inst
    t12_656 <= a31_516 when (SGT_i16_u1_652_wire(0) /=  '0') else a41_580;
    -- flow-through select operator MUX_663_inst
    out1_664 <= t11_648 when (SGT_i16_u1_660_wire(0) /=  '0') else t12_656;
    -- flow-through select operator MUX_671_inst
    t21_672 <= a12_392 when (SGT_i16_u1_668_wire(0) /=  '0') else a22_456;
    -- flow-through select operator MUX_679_inst
    t22_680 <= a32_520 when (SGT_i16_u1_676_wire(0) /=  '0') else a42_584;
    -- flow-through select operator MUX_687_inst
    out2_688 <= t21_672 when (SGT_i16_u1_684_wire(0) /=  '0') else t22_680;
    -- flow-through select operator MUX_695_inst
    t31_696 <= a13_396 when (SGT_i16_u1_692_wire(0) /=  '0') else a23_460;
    -- flow-through select operator MUX_703_inst
    t32_704 <= a33_524 when (SGT_i16_u1_700_wire(0) /=  '0') else a43_588;
    -- flow-through select operator MUX_711_inst
    out3_712 <= t31_696 when (SGT_i16_u1_708_wire(0) /=  '0') else t32_704;
    -- flow-through select operator MUX_719_inst
    t41_720 <= a14_400 when (SGT_i16_u1_716_wire(0) /=  '0') else a24_464;
    -- flow-through select operator MUX_727_inst
    t42_728 <= a34_528 when (SGT_i16_u1_724_wire(0) /=  '0') else a44_592;
    -- flow-through select operator MUX_735_inst
    out4_736 <= t41_720 when (SGT_i16_u1_732_wire(0) /=  '0') else t42_728;
    -- flow-through select operator MUX_743_inst
    t51_744 <= a15_404 when (SGT_i16_u1_740_wire(0) /=  '0') else a25_468;
    -- flow-through select operator MUX_751_inst
    t52_752 <= a35_532 when (SGT_i16_u1_748_wire(0) /=  '0') else a45_596;
    -- flow-through select operator MUX_759_inst
    out5_760 <= t51_744 when (SGT_i16_u1_756_wire(0) /=  '0') else t52_752;
    -- flow-through select operator MUX_767_inst
    t61_768 <= a16_408 when (SGT_i16_u1_764_wire(0) /=  '0') else a26_472;
    -- flow-through select operator MUX_775_inst
    t62_776 <= a36_536 when (SGT_i16_u1_772_wire(0) /=  '0') else a46_600;
    -- flow-through select operator MUX_783_inst
    out6_784 <= t61_768 when (SGT_i16_u1_780_wire(0) /=  '0') else t62_776;
    -- flow-through select operator MUX_791_inst
    t71_792 <= a17_412 when (SGT_i16_u1_788_wire(0) /=  '0') else a27_476;
    -- flow-through select operator MUX_799_inst
    t72_800 <= a37_540 when (SGT_i16_u1_796_wire(0) /=  '0') else a47_604;
    -- flow-through select operator MUX_807_inst
    out7_808 <= t71_792 when (SGT_i16_u1_804_wire(0) /=  '0') else t72_800;
    -- flow-through select operator MUX_815_inst
    t81_816 <= a18_416 when (SGT_i16_u1_812_wire(0) /=  '0') else a28_480;
    -- flow-through select operator MUX_823_inst
    t82_824 <= a38_544 when (SGT_i16_u1_820_wire(0) /=  '0') else a48_608;
    -- flow-through select operator MUX_831_inst
    out8_832 <= t81_816 when (SGT_i16_u1_828_wire(0) /=  '0') else t82_824;
    -- flow-through select operator MUX_839_inst
    t91_840 <= a19_420 when (SGT_i16_u1_836_wire(0) /=  '0') else a29_484;
    -- flow-through select operator MUX_847_inst
    t92_848 <= a39_548 when (SGT_i16_u1_844_wire(0) /=  '0') else a49_612;
    -- flow-through select operator MUX_855_inst
    out9_856 <= t91_840 when (SGT_i16_u1_852_wire(0) /=  '0') else t92_848;
    -- flow-through select operator MUX_863_inst
    t101_864 <= a110_424 when (SGT_i16_u1_860_wire(0) /=  '0') else a210_488;
    -- flow-through select operator MUX_871_inst
    t102_872 <= a310_552 when (SGT_i16_u1_868_wire(0) /=  '0') else a410_616;
    -- flow-through select operator MUX_879_inst
    out10_880 <= t101_864 when (SGT_i16_u1_876_wire(0) /=  '0') else t102_872;
    -- flow-through select operator MUX_887_inst
    t111_888 <= a111_428 when (SGT_i16_u1_884_wire(0) /=  '0') else a211_492;
    -- flow-through select operator MUX_895_inst
    t112_896 <= a311_556 when (SGT_i16_u1_892_wire(0) /=  '0') else a411_620;
    -- flow-through select operator MUX_903_inst
    out11_904 <= t111_888 when (SGT_i16_u1_900_wire(0) /=  '0') else t112_896;
    -- flow-through select operator MUX_911_inst
    t121_912 <= a112_432 when (SGT_i16_u1_908_wire(0) /=  '0') else a212_496;
    -- flow-through select operator MUX_919_inst
    t122_920 <= a312_560 when (SGT_i16_u1_916_wire(0) /=  '0') else a412_624;
    -- flow-through select operator MUX_927_inst
    out12_928 <= t121_912 when (SGT_i16_u1_924_wire(0) /=  '0') else t122_920;
    -- flow-through select operator MUX_935_inst
    t131_936 <= a113_436 when (SGT_i16_u1_932_wire(0) /=  '0') else a213_500;
    -- flow-through select operator MUX_943_inst
    t132_944 <= a313_564 when (SGT_i16_u1_940_wire(0) /=  '0') else a413_628;
    -- flow-through select operator MUX_951_inst
    out13_952 <= t131_936 when (SGT_i16_u1_948_wire(0) /=  '0') else t132_944;
    -- flow-through select operator MUX_959_inst
    t141_960 <= a114_440 when (SGT_i16_u1_956_wire(0) /=  '0') else a214_504;
    -- flow-through select operator MUX_967_inst
    t142_968 <= a314_568 when (SGT_i16_u1_964_wire(0) /=  '0') else a414_632;
    -- flow-through select operator MUX_975_inst
    out14_976 <= t141_960 when (SGT_i16_u1_972_wire(0) /=  '0') else t142_968;
    -- flow-through select operator MUX_983_inst
    t151_984 <= a115_444 when (SGT_i16_u1_980_wire(0) /=  '0') else a215_508;
    -- flow-through select operator MUX_991_inst
    t152_992 <= a315_572 when (SGT_i16_u1_988_wire(0) /=  '0') else a415_636;
    -- flow-through select operator MUX_999_inst
    out15_1000 <= t151_984 when (SGT_i16_u1_996_wire(0) /=  '0') else t152_992;
    slice_130_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_130_inst_req_0;
      slice_130_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_130_inst_req_1;
      slice_130_inst_ack_1<= update_ack(0);
      slice_130_inst: SliceSplitProtocol generic map(name => "slice_130_inst", in_data_width => 256, high_index => 255, low_index => 240, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_114, dout => sliced_v11_131, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_134_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_134_inst_req_0;
      slice_134_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_134_inst_req_1;
      slice_134_inst_ack_1<= update_ack(0);
      slice_134_inst: SliceSplitProtocol generic map(name => "slice_134_inst", in_data_width => 256, high_index => 239, low_index => 224, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_114, dout => sliced_v12_135, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_138_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_138_inst_req_0;
      slice_138_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_138_inst_req_1;
      slice_138_inst_ack_1<= update_ack(0);
      slice_138_inst: SliceSplitProtocol generic map(name => "slice_138_inst", in_data_width => 256, high_index => 223, low_index => 208, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_114, dout => sliced_v13_139, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_142_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_142_inst_req_0;
      slice_142_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_142_inst_req_1;
      slice_142_inst_ack_1<= update_ack(0);
      slice_142_inst: SliceSplitProtocol generic map(name => "slice_142_inst", in_data_width => 256, high_index => 207, low_index => 192, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_114, dout => sliced_v14_143, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_146_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_146_inst_req_0;
      slice_146_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_146_inst_req_1;
      slice_146_inst_ack_1<= update_ack(0);
      slice_146_inst: SliceSplitProtocol generic map(name => "slice_146_inst", in_data_width => 256, high_index => 191, low_index => 176, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_114, dout => sliced_v15_147, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_150_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_150_inst_req_0;
      slice_150_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_150_inst_req_1;
      slice_150_inst_ack_1<= update_ack(0);
      slice_150_inst: SliceSplitProtocol generic map(name => "slice_150_inst", in_data_width => 256, high_index => 175, low_index => 160, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_114, dout => sliced_v16_151, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_154_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_154_inst_req_0;
      slice_154_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_154_inst_req_1;
      slice_154_inst_ack_1<= update_ack(0);
      slice_154_inst: SliceSplitProtocol generic map(name => "slice_154_inst", in_data_width => 256, high_index => 159, low_index => 144, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_114, dout => sliced_v17_155, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_158_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_158_inst_req_0;
      slice_158_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_158_inst_req_1;
      slice_158_inst_ack_1<= update_ack(0);
      slice_158_inst: SliceSplitProtocol generic map(name => "slice_158_inst", in_data_width => 256, high_index => 143, low_index => 128, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_114, dout => sliced_v18_159, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_162_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_162_inst_req_0;
      slice_162_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_162_inst_req_1;
      slice_162_inst_ack_1<= update_ack(0);
      slice_162_inst: SliceSplitProtocol generic map(name => "slice_162_inst", in_data_width => 256, high_index => 127, low_index => 112, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_114, dout => sliced_v19_163, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_166_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_166_inst_req_0;
      slice_166_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_166_inst_req_1;
      slice_166_inst_ack_1<= update_ack(0);
      slice_166_inst: SliceSplitProtocol generic map(name => "slice_166_inst", in_data_width => 256, high_index => 111, low_index => 96, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_114, dout => sliced_v110_167, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_170_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_170_inst_req_0;
      slice_170_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_170_inst_req_1;
      slice_170_inst_ack_1<= update_ack(0);
      slice_170_inst: SliceSplitProtocol generic map(name => "slice_170_inst", in_data_width => 256, high_index => 95, low_index => 80, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_114, dout => sliced_v111_171, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_174_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_174_inst_req_0;
      slice_174_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_174_inst_req_1;
      slice_174_inst_ack_1<= update_ack(0);
      slice_174_inst: SliceSplitProtocol generic map(name => "slice_174_inst", in_data_width => 256, high_index => 79, low_index => 64, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_114, dout => sliced_v112_175, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_178_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_178_inst_req_0;
      slice_178_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_178_inst_req_1;
      slice_178_inst_ack_1<= update_ack(0);
      slice_178_inst: SliceSplitProtocol generic map(name => "slice_178_inst", in_data_width => 256, high_index => 63, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_114, dout => sliced_v113_179, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_182_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_182_inst_req_0;
      slice_182_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_182_inst_req_1;
      slice_182_inst_ack_1<= update_ack(0);
      slice_182_inst: SliceSplitProtocol generic map(name => "slice_182_inst", in_data_width => 256, high_index => 47, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_114, dout => sliced_v114_183, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_186_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_186_inst_req_0;
      slice_186_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_186_inst_req_1;
      slice_186_inst_ack_1<= update_ack(0);
      slice_186_inst: SliceSplitProtocol generic map(name => "slice_186_inst", in_data_width => 256, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_114, dout => sliced_v115_187, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_190_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_190_inst_req_0;
      slice_190_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_190_inst_req_1;
      slice_190_inst_ack_1<= update_ack(0);
      slice_190_inst: SliceSplitProtocol generic map(name => "slice_190_inst", in_data_width => 256, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_114, dout => sliced_v116_191, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_194_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_194_inst_req_0;
      slice_194_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_194_inst_req_1;
      slice_194_inst_ack_1<= update_ack(0);
      slice_194_inst: SliceSplitProtocol generic map(name => "slice_194_inst", in_data_width => 256, high_index => 255, low_index => 240, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_118, dout => sliced_v21_195, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_198_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_198_inst_req_0;
      slice_198_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_198_inst_req_1;
      slice_198_inst_ack_1<= update_ack(0);
      slice_198_inst: SliceSplitProtocol generic map(name => "slice_198_inst", in_data_width => 256, high_index => 239, low_index => 224, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_118, dout => sliced_v22_199, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_202_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_202_inst_req_0;
      slice_202_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_202_inst_req_1;
      slice_202_inst_ack_1<= update_ack(0);
      slice_202_inst: SliceSplitProtocol generic map(name => "slice_202_inst", in_data_width => 256, high_index => 223, low_index => 208, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_118, dout => sliced_v23_203, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_206_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_206_inst_req_0;
      slice_206_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_206_inst_req_1;
      slice_206_inst_ack_1<= update_ack(0);
      slice_206_inst: SliceSplitProtocol generic map(name => "slice_206_inst", in_data_width => 256, high_index => 207, low_index => 192, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_118, dout => sliced_v24_207, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_210_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_210_inst_req_0;
      slice_210_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_210_inst_req_1;
      slice_210_inst_ack_1<= update_ack(0);
      slice_210_inst: SliceSplitProtocol generic map(name => "slice_210_inst", in_data_width => 256, high_index => 191, low_index => 176, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_118, dout => sliced_v25_211, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_214_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_214_inst_req_0;
      slice_214_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_214_inst_req_1;
      slice_214_inst_ack_1<= update_ack(0);
      slice_214_inst: SliceSplitProtocol generic map(name => "slice_214_inst", in_data_width => 256, high_index => 175, low_index => 160, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_118, dout => sliced_v26_215, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_218_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_218_inst_req_0;
      slice_218_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_218_inst_req_1;
      slice_218_inst_ack_1<= update_ack(0);
      slice_218_inst: SliceSplitProtocol generic map(name => "slice_218_inst", in_data_width => 256, high_index => 159, low_index => 144, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_118, dout => sliced_v27_219, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_222_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_222_inst_req_0;
      slice_222_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_222_inst_req_1;
      slice_222_inst_ack_1<= update_ack(0);
      slice_222_inst: SliceSplitProtocol generic map(name => "slice_222_inst", in_data_width => 256, high_index => 143, low_index => 128, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_118, dout => sliced_v28_223, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_226_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_226_inst_req_0;
      slice_226_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_226_inst_req_1;
      slice_226_inst_ack_1<= update_ack(0);
      slice_226_inst: SliceSplitProtocol generic map(name => "slice_226_inst", in_data_width => 256, high_index => 127, low_index => 112, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_118, dout => sliced_v29_227, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_230_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_230_inst_req_0;
      slice_230_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_230_inst_req_1;
      slice_230_inst_ack_1<= update_ack(0);
      slice_230_inst: SliceSplitProtocol generic map(name => "slice_230_inst", in_data_width => 256, high_index => 111, low_index => 96, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_118, dout => sliced_v210_231, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_234_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_234_inst_req_0;
      slice_234_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_234_inst_req_1;
      slice_234_inst_ack_1<= update_ack(0);
      slice_234_inst: SliceSplitProtocol generic map(name => "slice_234_inst", in_data_width => 256, high_index => 95, low_index => 80, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_118, dout => sliced_v211_235, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_238_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_238_inst_req_0;
      slice_238_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_238_inst_req_1;
      slice_238_inst_ack_1<= update_ack(0);
      slice_238_inst: SliceSplitProtocol generic map(name => "slice_238_inst", in_data_width => 256, high_index => 79, low_index => 64, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_118, dout => sliced_v212_239, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_242_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_242_inst_req_0;
      slice_242_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_242_inst_req_1;
      slice_242_inst_ack_1<= update_ack(0);
      slice_242_inst: SliceSplitProtocol generic map(name => "slice_242_inst", in_data_width => 256, high_index => 63, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_118, dout => sliced_v213_243, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_246_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_246_inst_req_0;
      slice_246_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_246_inst_req_1;
      slice_246_inst_ack_1<= update_ack(0);
      slice_246_inst: SliceSplitProtocol generic map(name => "slice_246_inst", in_data_width => 256, high_index => 47, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_118, dout => sliced_v214_247, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_250_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_250_inst_req_0;
      slice_250_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_250_inst_req_1;
      slice_250_inst_ack_1<= update_ack(0);
      slice_250_inst: SliceSplitProtocol generic map(name => "slice_250_inst", in_data_width => 256, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_118, dout => sliced_v215_251, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_254_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_254_inst_req_0;
      slice_254_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_254_inst_req_1;
      slice_254_inst_ack_1<= update_ack(0);
      slice_254_inst: SliceSplitProtocol generic map(name => "slice_254_inst", in_data_width => 256, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_118, dout => sliced_v216_255, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_258_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_258_inst_req_0;
      slice_258_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_258_inst_req_1;
      slice_258_inst_ack_1<= update_ack(0);
      slice_258_inst: SliceSplitProtocol generic map(name => "slice_258_inst", in_data_width => 256, high_index => 255, low_index => 240, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_122, dout => sliced_v31_259, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_262_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_262_inst_req_0;
      slice_262_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_262_inst_req_1;
      slice_262_inst_ack_1<= update_ack(0);
      slice_262_inst: SliceSplitProtocol generic map(name => "slice_262_inst", in_data_width => 256, high_index => 239, low_index => 224, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_122, dout => sliced_v32_263, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_266_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_266_inst_req_0;
      slice_266_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_266_inst_req_1;
      slice_266_inst_ack_1<= update_ack(0);
      slice_266_inst: SliceSplitProtocol generic map(name => "slice_266_inst", in_data_width => 256, high_index => 223, low_index => 208, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_122, dout => sliced_v33_267, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_270_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_270_inst_req_0;
      slice_270_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_270_inst_req_1;
      slice_270_inst_ack_1<= update_ack(0);
      slice_270_inst: SliceSplitProtocol generic map(name => "slice_270_inst", in_data_width => 256, high_index => 207, low_index => 192, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_122, dout => sliced_v34_271, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_274_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_274_inst_req_0;
      slice_274_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_274_inst_req_1;
      slice_274_inst_ack_1<= update_ack(0);
      slice_274_inst: SliceSplitProtocol generic map(name => "slice_274_inst", in_data_width => 256, high_index => 191, low_index => 176, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_122, dout => sliced_v35_275, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_278_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_278_inst_req_0;
      slice_278_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_278_inst_req_1;
      slice_278_inst_ack_1<= update_ack(0);
      slice_278_inst: SliceSplitProtocol generic map(name => "slice_278_inst", in_data_width => 256, high_index => 175, low_index => 160, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_122, dout => sliced_v36_279, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_282_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_282_inst_req_0;
      slice_282_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_282_inst_req_1;
      slice_282_inst_ack_1<= update_ack(0);
      slice_282_inst: SliceSplitProtocol generic map(name => "slice_282_inst", in_data_width => 256, high_index => 159, low_index => 144, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_122, dout => sliced_v37_283, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_286_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_286_inst_req_0;
      slice_286_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_286_inst_req_1;
      slice_286_inst_ack_1<= update_ack(0);
      slice_286_inst: SliceSplitProtocol generic map(name => "slice_286_inst", in_data_width => 256, high_index => 143, low_index => 128, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_122, dout => sliced_v38_287, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_290_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_290_inst_req_0;
      slice_290_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_290_inst_req_1;
      slice_290_inst_ack_1<= update_ack(0);
      slice_290_inst: SliceSplitProtocol generic map(name => "slice_290_inst", in_data_width => 256, high_index => 127, low_index => 112, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_122, dout => sliced_v39_291, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_294_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_294_inst_req_0;
      slice_294_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_294_inst_req_1;
      slice_294_inst_ack_1<= update_ack(0);
      slice_294_inst: SliceSplitProtocol generic map(name => "slice_294_inst", in_data_width => 256, high_index => 111, low_index => 96, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_122, dout => sliced_v310_295, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_298_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_298_inst_req_0;
      slice_298_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_298_inst_req_1;
      slice_298_inst_ack_1<= update_ack(0);
      slice_298_inst: SliceSplitProtocol generic map(name => "slice_298_inst", in_data_width => 256, high_index => 95, low_index => 80, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_122, dout => sliced_v311_299, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_302_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_302_inst_req_0;
      slice_302_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_302_inst_req_1;
      slice_302_inst_ack_1<= update_ack(0);
      slice_302_inst: SliceSplitProtocol generic map(name => "slice_302_inst", in_data_width => 256, high_index => 79, low_index => 64, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_122, dout => sliced_v312_303, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_306_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_306_inst_req_0;
      slice_306_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_306_inst_req_1;
      slice_306_inst_ack_1<= update_ack(0);
      slice_306_inst: SliceSplitProtocol generic map(name => "slice_306_inst", in_data_width => 256, high_index => 63, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_122, dout => sliced_v313_307, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_310_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_310_inst_req_0;
      slice_310_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_310_inst_req_1;
      slice_310_inst_ack_1<= update_ack(0);
      slice_310_inst: SliceSplitProtocol generic map(name => "slice_310_inst", in_data_width => 256, high_index => 47, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_122, dout => sliced_v314_311, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_314_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_314_inst_req_0;
      slice_314_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_314_inst_req_1;
      slice_314_inst_ack_1<= update_ack(0);
      slice_314_inst: SliceSplitProtocol generic map(name => "slice_314_inst", in_data_width => 256, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_122, dout => sliced_v315_315, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_318_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_318_inst_req_0;
      slice_318_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_318_inst_req_1;
      slice_318_inst_ack_1<= update_ack(0);
      slice_318_inst: SliceSplitProtocol generic map(name => "slice_318_inst", in_data_width => 256, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_122, dout => sliced_v316_319, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_322_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_322_inst_req_0;
      slice_322_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_322_inst_req_1;
      slice_322_inst_ack_1<= update_ack(0);
      slice_322_inst: SliceSplitProtocol generic map(name => "slice_322_inst", in_data_width => 256, high_index => 255, low_index => 240, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_126, dout => sliced_v41_323, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_326_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_326_inst_req_0;
      slice_326_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_326_inst_req_1;
      slice_326_inst_ack_1<= update_ack(0);
      slice_326_inst: SliceSplitProtocol generic map(name => "slice_326_inst", in_data_width => 256, high_index => 239, low_index => 224, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_126, dout => sliced_v42_327, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_330_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_330_inst_req_0;
      slice_330_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_330_inst_req_1;
      slice_330_inst_ack_1<= update_ack(0);
      slice_330_inst: SliceSplitProtocol generic map(name => "slice_330_inst", in_data_width => 256, high_index => 223, low_index => 208, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_126, dout => sliced_v43_331, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_334_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_334_inst_req_0;
      slice_334_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_334_inst_req_1;
      slice_334_inst_ack_1<= update_ack(0);
      slice_334_inst: SliceSplitProtocol generic map(name => "slice_334_inst", in_data_width => 256, high_index => 207, low_index => 192, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_126, dout => sliced_v44_335, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_338_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_338_inst_req_0;
      slice_338_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_338_inst_req_1;
      slice_338_inst_ack_1<= update_ack(0);
      slice_338_inst: SliceSplitProtocol generic map(name => "slice_338_inst", in_data_width => 256, high_index => 191, low_index => 176, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_126, dout => sliced_v45_339, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_342_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_342_inst_req_0;
      slice_342_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_342_inst_req_1;
      slice_342_inst_ack_1<= update_ack(0);
      slice_342_inst: SliceSplitProtocol generic map(name => "slice_342_inst", in_data_width => 256, high_index => 175, low_index => 160, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_126, dout => sliced_v46_343, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_346_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_346_inst_req_0;
      slice_346_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_346_inst_req_1;
      slice_346_inst_ack_1<= update_ack(0);
      slice_346_inst: SliceSplitProtocol generic map(name => "slice_346_inst", in_data_width => 256, high_index => 159, low_index => 144, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_126, dout => sliced_v47_347, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_350_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_350_inst_req_0;
      slice_350_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_350_inst_req_1;
      slice_350_inst_ack_1<= update_ack(0);
      slice_350_inst: SliceSplitProtocol generic map(name => "slice_350_inst", in_data_width => 256, high_index => 143, low_index => 128, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_126, dout => sliced_v48_351, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_354_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_354_inst_req_0;
      slice_354_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_354_inst_req_1;
      slice_354_inst_ack_1<= update_ack(0);
      slice_354_inst: SliceSplitProtocol generic map(name => "slice_354_inst", in_data_width => 256, high_index => 127, low_index => 112, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_126, dout => sliced_v49_355, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_358_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_358_inst_req_0;
      slice_358_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_358_inst_req_1;
      slice_358_inst_ack_1<= update_ack(0);
      slice_358_inst: SliceSplitProtocol generic map(name => "slice_358_inst", in_data_width => 256, high_index => 111, low_index => 96, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_126, dout => sliced_v410_359, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_362_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_362_inst_req_0;
      slice_362_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_362_inst_req_1;
      slice_362_inst_ack_1<= update_ack(0);
      slice_362_inst: SliceSplitProtocol generic map(name => "slice_362_inst", in_data_width => 256, high_index => 95, low_index => 80, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_126, dout => sliced_v411_363, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_366_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_366_inst_req_0;
      slice_366_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_366_inst_req_1;
      slice_366_inst_ack_1<= update_ack(0);
      slice_366_inst: SliceSplitProtocol generic map(name => "slice_366_inst", in_data_width => 256, high_index => 79, low_index => 64, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_126, dout => sliced_v412_367, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_370_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_370_inst_req_0;
      slice_370_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_370_inst_req_1;
      slice_370_inst_ack_1<= update_ack(0);
      slice_370_inst: SliceSplitProtocol generic map(name => "slice_370_inst", in_data_width => 256, high_index => 63, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_126, dout => sliced_v413_371, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_374_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_374_inst_req_0;
      slice_374_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_374_inst_req_1;
      slice_374_inst_ack_1<= update_ack(0);
      slice_374_inst: SliceSplitProtocol generic map(name => "slice_374_inst", in_data_width => 256, high_index => 47, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_126, dout => sliced_v414_375, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_378_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_378_inst_req_0;
      slice_378_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_378_inst_req_1;
      slice_378_inst_ack_1<= update_ack(0);
      slice_378_inst: SliceSplitProtocol generic map(name => "slice_378_inst", in_data_width => 256, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_126, dout => sliced_v415_379, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_382_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_382_inst_req_0;
      slice_382_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_382_inst_req_1;
      slice_382_inst_ack_1<= update_ack(0);
      slice_382_inst: SliceSplitProtocol generic map(name => "slice_382_inst", in_data_width => 256, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_126, dout => sliced_v416_383, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    W_myptr5_1032_delayed_8_0_1032_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_myptr5_1032_delayed_8_0_1032_inst_req_0;
      W_myptr5_1032_delayed_8_0_1032_inst_ack_0<= wack(0);
      rreq(0) <= W_myptr5_1032_delayed_8_0_1032_inst_req_1;
      W_myptr5_1032_delayed_8_0_1032_inst_ack_1<= rack(0);
      W_myptr5_1032_delayed_8_0_1032_inst : InterlockBuffer generic map ( -- 
        name => "W_myptr5_1032_delayed_8_0_1032_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => myptr5_1031,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr5_1032_delayed_8_0_1034,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_myptr6_1055_delayed_8_0_1058_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_myptr6_1055_delayed_8_0_1058_inst_req_0;
      W_myptr6_1055_delayed_8_0_1058_inst_ack_0<= wack(0);
      rreq(0) <= W_myptr6_1055_delayed_8_0_1058_inst_req_1;
      W_myptr6_1055_delayed_8_0_1058_inst_ack_1<= rack(0);
      W_myptr6_1055_delayed_8_0_1058_inst : InterlockBuffer generic map ( -- 
        name => "W_myptr6_1055_delayed_8_0_1058_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => myptr6_1057,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr6_1055_delayed_8_0_1060,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_myptr7_1078_delayed_8_0_1084_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_myptr7_1078_delayed_8_0_1084_inst_req_0;
      W_myptr7_1078_delayed_8_0_1084_inst_ack_0<= wack(0);
      rreq(0) <= W_myptr7_1078_delayed_8_0_1084_inst_req_1;
      W_myptr7_1078_delayed_8_0_1084_inst_ack_1<= rack(0);
      W_myptr7_1078_delayed_8_0_1084_inst : InterlockBuffer generic map ( -- 
        name => "W_myptr7_1078_delayed_8_0_1084_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => myptr7_1083,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr7_1078_delayed_8_0_1086,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_myptr8_1101_delayed_8_0_1110_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_myptr8_1101_delayed_8_0_1110_inst_req_0;
      W_myptr8_1101_delayed_8_0_1110_inst_ack_0<= wack(0);
      rreq(0) <= W_myptr8_1101_delayed_8_0_1110_inst_req_1;
      W_myptr8_1101_delayed_8_0_1110_inst_ack_1<= rack(0);
      W_myptr8_1101_delayed_8_0_1110_inst : InterlockBuffer generic map ( -- 
        name => "W_myptr8_1101_delayed_8_0_1110_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => myptr8_1109,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr8_1101_delayed_8_0_1112,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_102_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_102_final_reg_req_0;
      addr_of_102_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_102_final_reg_req_1;
      addr_of_102_final_reg_ack_1<= rack(0);
      addr_of_102_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_102_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_101_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr3_103,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1030_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1030_final_reg_req_0;
      addr_of_1030_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1030_final_reg_req_1;
      addr_of_1030_final_reg_ack_1<= rack(0);
      addr_of_1030_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1030_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1029_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr5_1031,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1056_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1056_final_reg_req_0;
      addr_of_1056_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1056_final_reg_req_1;
      addr_of_1056_final_reg_ack_1<= rack(0);
      addr_of_1056_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1056_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1055_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr6_1057,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1082_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1082_final_reg_req_0;
      addr_of_1082_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1082_final_reg_req_1;
      addr_of_1082_final_reg_ack_1<= rack(0);
      addr_of_1082_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1082_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1081_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr7_1083,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_109_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_109_final_reg_req_0;
      addr_of_109_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_109_final_reg_req_1;
      addr_of_109_final_reg_ack_1<= rack(0);
      addr_of_109_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_109_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_108_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr4_110,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1108_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1108_final_reg_req_0;
      addr_of_1108_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1108_final_reg_req_1;
      addr_of_1108_final_reg_ack_1<= rack(0);
      addr_of_1108_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1108_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1107_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr8_1109,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_88_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_88_final_reg_req_0;
      addr_of_88_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_88_final_reg_req_1;
      addr_of_88_final_reg_ack_1<= rack(0);
      addr_of_88_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_88_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_87_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr1_89,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_95_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_95_final_reg_req_0;
      addr_of_95_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_95_final_reg_req_1;
      addr_of_95_final_reg_ack_1<= rack(0);
      addr_of_95_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_95_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_94_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr2_96,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1038_inst
    process(out1_664) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out1_664(15 downto 0);
      type_cast_1038_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1040_inst
    process(out2_688) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out2_688(15 downto 0);
      type_cast_1040_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1043_inst
    process(out3_712) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out3_712(15 downto 0);
      type_cast_1043_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1045_inst
    process(out4_736) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out4_736(15 downto 0);
      type_cast_1045_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1064_inst
    process(out5_760) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out5_760(15 downto 0);
      type_cast_1064_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1066_inst
    process(out6_784) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out6_784(15 downto 0);
      type_cast_1066_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1069_inst
    process(out7_808) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out7_808(15 downto 0);
      type_cast_1069_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1071_inst
    process(out8_832) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out8_832(15 downto 0);
      type_cast_1071_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1090_inst
    process(out9_856) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out9_856(15 downto 0);
      type_cast_1090_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1092_inst
    process(out10_880) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out10_880(15 downto 0);
      type_cast_1092_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1095_inst
    process(out11_904) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out11_904(15 downto 0);
      type_cast_1095_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1097_inst
    process(out12_928) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out12_928(15 downto 0);
      type_cast_1097_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1116_inst
    process(out13_952) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out13_952(15 downto 0);
      type_cast_1116_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1118_inst
    process(out14_976) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out14_976(15 downto 0);
      type_cast_1118_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1121_inst
    process(out15_1000) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out15_1000(15 downto 0);
      type_cast_1121_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1123_inst
    process(out16_1024) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out16_1024(15 downto 0);
      type_cast_1123_wire <= tmp_var; -- 
    end process;
    type_cast_1129_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1129_inst_req_0;
      type_cast_1129_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1129_inst_req_1;
      type_cast_1129_inst_ack_1<= rack(0);
      type_cast_1129_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1129_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => out1_664,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_buffer,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_387_inst
    process(sliced_v11_131) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v11_131(15 downto 0);
      a11_388 <= tmp_var; -- 
    end process;
    -- interlock type_cast_391_inst
    process(sliced_v12_135) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v12_135(15 downto 0);
      a12_392 <= tmp_var; -- 
    end process;
    -- interlock type_cast_395_inst
    process(sliced_v13_139) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v13_139(15 downto 0);
      a13_396 <= tmp_var; -- 
    end process;
    -- interlock type_cast_399_inst
    process(sliced_v14_143) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v14_143(15 downto 0);
      a14_400 <= tmp_var; -- 
    end process;
    -- interlock type_cast_403_inst
    process(sliced_v15_147) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v15_147(15 downto 0);
      a15_404 <= tmp_var; -- 
    end process;
    -- interlock type_cast_407_inst
    process(sliced_v16_151) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v16_151(15 downto 0);
      a16_408 <= tmp_var; -- 
    end process;
    -- interlock type_cast_411_inst
    process(sliced_v17_155) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v17_155(15 downto 0);
      a17_412 <= tmp_var; -- 
    end process;
    -- interlock type_cast_415_inst
    process(sliced_v18_159) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v18_159(15 downto 0);
      a18_416 <= tmp_var; -- 
    end process;
    -- interlock type_cast_419_inst
    process(sliced_v19_163) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v19_163(15 downto 0);
      a19_420 <= tmp_var; -- 
    end process;
    -- interlock type_cast_423_inst
    process(sliced_v110_167) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v110_167(15 downto 0);
      a110_424 <= tmp_var; -- 
    end process;
    -- interlock type_cast_427_inst
    process(sliced_v111_171) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v111_171(15 downto 0);
      a111_428 <= tmp_var; -- 
    end process;
    -- interlock type_cast_431_inst
    process(sliced_v112_175) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v112_175(15 downto 0);
      a112_432 <= tmp_var; -- 
    end process;
    -- interlock type_cast_435_inst
    process(sliced_v113_179) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v113_179(15 downto 0);
      a113_436 <= tmp_var; -- 
    end process;
    -- interlock type_cast_439_inst
    process(sliced_v114_183) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v114_183(15 downto 0);
      a114_440 <= tmp_var; -- 
    end process;
    -- interlock type_cast_443_inst
    process(sliced_v115_187) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v115_187(15 downto 0);
      a115_444 <= tmp_var; -- 
    end process;
    -- interlock type_cast_447_inst
    process(sliced_v116_191) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v116_191(15 downto 0);
      a116_448 <= tmp_var; -- 
    end process;
    -- interlock type_cast_451_inst
    process(sliced_v21_195) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v21_195(15 downto 0);
      a21_452 <= tmp_var; -- 
    end process;
    -- interlock type_cast_455_inst
    process(sliced_v22_199) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v22_199(15 downto 0);
      a22_456 <= tmp_var; -- 
    end process;
    -- interlock type_cast_459_inst
    process(sliced_v23_203) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v23_203(15 downto 0);
      a23_460 <= tmp_var; -- 
    end process;
    -- interlock type_cast_463_inst
    process(sliced_v24_207) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v24_207(15 downto 0);
      a24_464 <= tmp_var; -- 
    end process;
    -- interlock type_cast_467_inst
    process(sliced_v25_211) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v25_211(15 downto 0);
      a25_468 <= tmp_var; -- 
    end process;
    -- interlock type_cast_471_inst
    process(sliced_v26_215) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v26_215(15 downto 0);
      a26_472 <= tmp_var; -- 
    end process;
    -- interlock type_cast_475_inst
    process(sliced_v27_219) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v27_219(15 downto 0);
      a27_476 <= tmp_var; -- 
    end process;
    -- interlock type_cast_479_inst
    process(sliced_v28_223) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v28_223(15 downto 0);
      a28_480 <= tmp_var; -- 
    end process;
    -- interlock type_cast_483_inst
    process(sliced_v29_227) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v29_227(15 downto 0);
      a29_484 <= tmp_var; -- 
    end process;
    -- interlock type_cast_487_inst
    process(sliced_v210_231) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v210_231(15 downto 0);
      a210_488 <= tmp_var; -- 
    end process;
    -- interlock type_cast_491_inst
    process(sliced_v211_235) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v211_235(15 downto 0);
      a211_492 <= tmp_var; -- 
    end process;
    -- interlock type_cast_495_inst
    process(sliced_v212_239) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v212_239(15 downto 0);
      a212_496 <= tmp_var; -- 
    end process;
    -- interlock type_cast_499_inst
    process(sliced_v213_243) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v213_243(15 downto 0);
      a213_500 <= tmp_var; -- 
    end process;
    -- interlock type_cast_503_inst
    process(sliced_v214_247) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v214_247(15 downto 0);
      a214_504 <= tmp_var; -- 
    end process;
    -- interlock type_cast_507_inst
    process(sliced_v215_251) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v215_251(15 downto 0);
      a215_508 <= tmp_var; -- 
    end process;
    -- interlock type_cast_511_inst
    process(sliced_v216_255) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v216_255(15 downto 0);
      a216_512 <= tmp_var; -- 
    end process;
    -- interlock type_cast_515_inst
    process(sliced_v31_259) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v31_259(15 downto 0);
      a31_516 <= tmp_var; -- 
    end process;
    -- interlock type_cast_519_inst
    process(sliced_v32_263) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v32_263(15 downto 0);
      a32_520 <= tmp_var; -- 
    end process;
    -- interlock type_cast_523_inst
    process(sliced_v33_267) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v33_267(15 downto 0);
      a33_524 <= tmp_var; -- 
    end process;
    -- interlock type_cast_527_inst
    process(sliced_v34_271) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v34_271(15 downto 0);
      a34_528 <= tmp_var; -- 
    end process;
    -- interlock type_cast_531_inst
    process(sliced_v35_275) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v35_275(15 downto 0);
      a35_532 <= tmp_var; -- 
    end process;
    -- interlock type_cast_535_inst
    process(sliced_v36_279) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v36_279(15 downto 0);
      a36_536 <= tmp_var; -- 
    end process;
    -- interlock type_cast_539_inst
    process(sliced_v37_283) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v37_283(15 downto 0);
      a37_540 <= tmp_var; -- 
    end process;
    -- interlock type_cast_543_inst
    process(sliced_v38_287) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v38_287(15 downto 0);
      a38_544 <= tmp_var; -- 
    end process;
    -- interlock type_cast_547_inst
    process(sliced_v39_291) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v39_291(15 downto 0);
      a39_548 <= tmp_var; -- 
    end process;
    -- interlock type_cast_551_inst
    process(sliced_v310_295) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v310_295(15 downto 0);
      a310_552 <= tmp_var; -- 
    end process;
    -- interlock type_cast_555_inst
    process(sliced_v311_299) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v311_299(15 downto 0);
      a311_556 <= tmp_var; -- 
    end process;
    -- interlock type_cast_559_inst
    process(sliced_v312_303) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v312_303(15 downto 0);
      a312_560 <= tmp_var; -- 
    end process;
    -- interlock type_cast_563_inst
    process(sliced_v313_307) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v313_307(15 downto 0);
      a313_564 <= tmp_var; -- 
    end process;
    -- interlock type_cast_567_inst
    process(sliced_v314_311) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v314_311(15 downto 0);
      a314_568 <= tmp_var; -- 
    end process;
    -- interlock type_cast_571_inst
    process(sliced_v315_315) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v315_315(15 downto 0);
      a315_572 <= tmp_var; -- 
    end process;
    -- interlock type_cast_575_inst
    process(sliced_v316_319) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v316_319(15 downto 0);
      a316_576 <= tmp_var; -- 
    end process;
    -- interlock type_cast_579_inst
    process(sliced_v41_323) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v41_323(15 downto 0);
      a41_580 <= tmp_var; -- 
    end process;
    -- interlock type_cast_583_inst
    process(sliced_v42_327) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v42_327(15 downto 0);
      a42_584 <= tmp_var; -- 
    end process;
    -- interlock type_cast_587_inst
    process(sliced_v43_331) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v43_331(15 downto 0);
      a43_588 <= tmp_var; -- 
    end process;
    -- interlock type_cast_591_inst
    process(sliced_v44_335) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v44_335(15 downto 0);
      a44_592 <= tmp_var; -- 
    end process;
    -- interlock type_cast_595_inst
    process(sliced_v45_339) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v45_339(15 downto 0);
      a45_596 <= tmp_var; -- 
    end process;
    -- interlock type_cast_599_inst
    process(sliced_v46_343) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v46_343(15 downto 0);
      a46_600 <= tmp_var; -- 
    end process;
    -- interlock type_cast_603_inst
    process(sliced_v47_347) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v47_347(15 downto 0);
      a47_604 <= tmp_var; -- 
    end process;
    -- interlock type_cast_607_inst
    process(sliced_v48_351) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v48_351(15 downto 0);
      a48_608 <= tmp_var; -- 
    end process;
    -- interlock type_cast_611_inst
    process(sliced_v49_355) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v49_355(15 downto 0);
      a49_612 <= tmp_var; -- 
    end process;
    -- interlock type_cast_615_inst
    process(sliced_v410_359) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v410_359(15 downto 0);
      a410_616 <= tmp_var; -- 
    end process;
    -- interlock type_cast_619_inst
    process(sliced_v411_363) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v411_363(15 downto 0);
      a411_620 <= tmp_var; -- 
    end process;
    -- interlock type_cast_623_inst
    process(sliced_v412_367) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v412_367(15 downto 0);
      a412_624 <= tmp_var; -- 
    end process;
    -- interlock type_cast_627_inst
    process(sliced_v413_371) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v413_371(15 downto 0);
      a413_628 <= tmp_var; -- 
    end process;
    -- interlock type_cast_631_inst
    process(sliced_v414_375) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v414_375(15 downto 0);
      a414_632 <= tmp_var; -- 
    end process;
    -- interlock type_cast_635_inst
    process(sliced_v415_379) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v415_379(15 downto 0);
      a415_636 <= tmp_var; -- 
    end process;
    -- interlock type_cast_639_inst
    process(sliced_v416_383) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v416_383(15 downto 0);
      a416_640 <= tmp_var; -- 
    end process;
    -- equivalence array_obj_ref_101_index_1_rename
    process(R_addr3_100_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr3_100_resized;
      ov(13 downto 0) := iv;
      R_addr3_100_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_101_index_1_resize
    process(addr3_buffer) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr3_buffer;
      ov := iv(13 downto 0);
      R_addr3_100_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_101_root_address_inst
    process(array_obj_ref_101_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_101_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_101_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1029_index_1_rename
    process(R_addr_1028_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr_1028_resized;
      ov(13 downto 0) := iv;
      R_addr_1028_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1029_index_1_resize
    process(addr_buffer) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr_buffer;
      ov := iv(13 downto 0);
      R_addr_1028_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1029_root_address_inst
    process(array_obj_ref_1029_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1029_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1029_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1055_index_1_rename
    process(ADD_u32_u32_1054_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ADD_u32_u32_1054_resized;
      ov(13 downto 0) := iv;
      ADD_u32_u32_1054_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1055_index_1_resize
    process(ADD_u32_u32_1054_wire) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ADD_u32_u32_1054_wire;
      ov := iv(13 downto 0);
      ADD_u32_u32_1054_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1055_root_address_inst
    process(array_obj_ref_1055_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1055_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1055_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1081_index_1_rename
    process(ADD_u32_u32_1080_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ADD_u32_u32_1080_resized;
      ov(13 downto 0) := iv;
      ADD_u32_u32_1080_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1081_index_1_resize
    process(ADD_u32_u32_1080_wire) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ADD_u32_u32_1080_wire;
      ov := iv(13 downto 0);
      ADD_u32_u32_1080_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1081_root_address_inst
    process(array_obj_ref_1081_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1081_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1081_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_108_index_1_rename
    process(R_addr4_107_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr4_107_resized;
      ov(13 downto 0) := iv;
      R_addr4_107_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_108_index_1_resize
    process(addr4_buffer) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr4_buffer;
      ov := iv(13 downto 0);
      R_addr4_107_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_108_root_address_inst
    process(array_obj_ref_108_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_108_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_108_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1107_index_1_rename
    process(ADD_u32_u32_1106_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ADD_u32_u32_1106_resized;
      ov(13 downto 0) := iv;
      ADD_u32_u32_1106_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1107_index_1_resize
    process(ADD_u32_u32_1106_wire) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ADD_u32_u32_1106_wire;
      ov := iv(13 downto 0);
      ADD_u32_u32_1106_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1107_root_address_inst
    process(array_obj_ref_1107_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1107_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1107_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_87_index_1_rename
    process(R_addr1_86_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr1_86_resized;
      ov(13 downto 0) := iv;
      R_addr1_86_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_87_index_1_resize
    process(addr1_buffer) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr1_buffer;
      ov := iv(13 downto 0);
      R_addr1_86_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_87_root_address_inst
    process(array_obj_ref_87_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_87_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_87_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_94_index_1_rename
    process(R_addr2_93_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr2_93_resized;
      ov(13 downto 0) := iv;
      R_addr2_93_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_94_index_1_resize
    process(addr2_buffer) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr2_buffer;
      ov := iv(13 downto 0);
      R_addr2_93_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_94_root_address_inst
    process(array_obj_ref_94_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_94_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_94_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1036_addr_0
    process(ptr_deref_1036_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1036_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1036_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1036_base_resize
    process(myptr5_1032_delayed_8_0_1034) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := myptr5_1032_delayed_8_0_1034;
      ov := iv(13 downto 0);
      ptr_deref_1036_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1036_gather_scatter
    process(CONCAT_u32_u64_1047_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := CONCAT_u32_u64_1047_wire;
      ov(63 downto 0) := iv;
      ptr_deref_1036_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1036_root_address_inst
    process(ptr_deref_1036_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1036_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1036_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1062_addr_0
    process(ptr_deref_1062_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1062_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1062_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1062_base_resize
    process(myptr6_1055_delayed_8_0_1060) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := myptr6_1055_delayed_8_0_1060;
      ov := iv(13 downto 0);
      ptr_deref_1062_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1062_gather_scatter
    process(CONCAT_u32_u64_1073_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := CONCAT_u32_u64_1073_wire;
      ov(63 downto 0) := iv;
      ptr_deref_1062_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1062_root_address_inst
    process(ptr_deref_1062_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1062_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1062_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1088_addr_0
    process(ptr_deref_1088_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1088_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1088_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1088_base_resize
    process(myptr7_1078_delayed_8_0_1086) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := myptr7_1078_delayed_8_0_1086;
      ov := iv(13 downto 0);
      ptr_deref_1088_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1088_gather_scatter
    process(CONCAT_u32_u64_1099_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := CONCAT_u32_u64_1099_wire;
      ov(63 downto 0) := iv;
      ptr_deref_1088_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1088_root_address_inst
    process(ptr_deref_1088_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1088_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1088_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1114_addr_0
    process(ptr_deref_1114_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1114_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1114_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1114_base_resize
    process(myptr8_1101_delayed_8_0_1112) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := myptr8_1101_delayed_8_0_1112;
      ov := iv(13 downto 0);
      ptr_deref_1114_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1114_gather_scatter
    process(CONCAT_u32_u64_1125_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := CONCAT_u32_u64_1125_wire;
      ov(63 downto 0) := iv;
      ptr_deref_1114_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1114_root_address_inst
    process(ptr_deref_1114_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1114_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1114_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_113_addr_0
    process(ptr_deref_113_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_113_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_113_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_113_base_resize
    process(myptr1_89) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := myptr1_89;
      ov := iv(13 downto 0);
      ptr_deref_113_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_113_gather_scatter
    process(ptr_deref_113_data_0) --
      variable iv : std_logic_vector(255 downto 0);
      variable ov : std_logic_vector(255 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_113_data_0;
      ov(255 downto 0) := iv;
      c1_114 <= ov(255 downto 0);
      --
    end process;
    -- equivalence ptr_deref_113_root_address_inst
    process(ptr_deref_113_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_113_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_113_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_117_addr_0
    process(ptr_deref_117_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_117_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_117_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_117_base_resize
    process(myptr2_96) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := myptr2_96;
      ov := iv(13 downto 0);
      ptr_deref_117_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_117_gather_scatter
    process(ptr_deref_117_data_0) --
      variable iv : std_logic_vector(255 downto 0);
      variable ov : std_logic_vector(255 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_117_data_0;
      ov(255 downto 0) := iv;
      c2_118 <= ov(255 downto 0);
      --
    end process;
    -- equivalence ptr_deref_117_root_address_inst
    process(ptr_deref_117_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_117_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_117_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_121_addr_0
    process(ptr_deref_121_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_121_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_121_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_121_base_resize
    process(myptr3_103) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := myptr3_103;
      ov := iv(13 downto 0);
      ptr_deref_121_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_121_gather_scatter
    process(ptr_deref_121_data_0) --
      variable iv : std_logic_vector(255 downto 0);
      variable ov : std_logic_vector(255 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_121_data_0;
      ov(255 downto 0) := iv;
      c3_122 <= ov(255 downto 0);
      --
    end process;
    -- equivalence ptr_deref_121_root_address_inst
    process(ptr_deref_121_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_121_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_121_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_125_addr_0
    process(ptr_deref_125_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_125_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_125_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_125_base_resize
    process(myptr4_110) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := myptr4_110;
      ov := iv(13 downto 0);
      ptr_deref_125_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_125_gather_scatter
    process(ptr_deref_125_data_0) --
      variable iv : std_logic_vector(255 downto 0);
      variable ov : std_logic_vector(255 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_125_data_0;
      ov(255 downto 0) := iv;
      c4_126 <= ov(255 downto 0);
      --
    end process;
    -- equivalence ptr_deref_125_root_address_inst
    process(ptr_deref_125_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_125_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_125_root_address <= ov(13 downto 0);
      --
    end process;
    -- binary operator ADD_u32_u32_1054_inst
    process(addr_buffer) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(addr_buffer, konst_1053_wire_constant, tmp_var);
      ADD_u32_u32_1054_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1080_inst
    process(addr_buffer) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(addr_buffer, konst_1079_wire_constant, tmp_var);
      ADD_u32_u32_1080_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1106_inst
    process(addr_buffer) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(addr_buffer, konst_1105_wire_constant, tmp_var);
      ADD_u32_u32_1106_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_1041_inst
    process(type_cast_1038_wire, type_cast_1040_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1038_wire, type_cast_1040_wire, tmp_var);
      CONCAT_u16_u32_1041_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_1046_inst
    process(type_cast_1043_wire, type_cast_1045_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1043_wire, type_cast_1045_wire, tmp_var);
      CONCAT_u16_u32_1046_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_1067_inst
    process(type_cast_1064_wire, type_cast_1066_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1064_wire, type_cast_1066_wire, tmp_var);
      CONCAT_u16_u32_1067_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_1072_inst
    process(type_cast_1069_wire, type_cast_1071_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1069_wire, type_cast_1071_wire, tmp_var);
      CONCAT_u16_u32_1072_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_1093_inst
    process(type_cast_1090_wire, type_cast_1092_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1090_wire, type_cast_1092_wire, tmp_var);
      CONCAT_u16_u32_1093_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_1098_inst
    process(type_cast_1095_wire, type_cast_1097_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1095_wire, type_cast_1097_wire, tmp_var);
      CONCAT_u16_u32_1098_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_1119_inst
    process(type_cast_1116_wire, type_cast_1118_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1116_wire, type_cast_1118_wire, tmp_var);
      CONCAT_u16_u32_1119_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_1124_inst
    process(type_cast_1121_wire, type_cast_1123_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1121_wire, type_cast_1123_wire, tmp_var);
      CONCAT_u16_u32_1124_wire <= tmp_var; --
    end process;
    -- shared split operator group (11) : CONCAT_u32_u64_1047_inst 
    ApConcat_group_11: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u16_u32_1041_wire & CONCAT_u16_u32_1046_wire;
      CONCAT_u32_u64_1047_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u32_u64_1047_inst_req_0;
      CONCAT_u32_u64_1047_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u32_u64_1047_inst_req_1;
      CONCAT_u32_u64_1047_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_11_gI: SplitGuardInterface generic map(name => "ApConcat_group_11_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_11",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared split operator group (12) : CONCAT_u32_u64_1073_inst 
    ApConcat_group_12: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u16_u32_1067_wire & CONCAT_u16_u32_1072_wire;
      CONCAT_u32_u64_1073_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u32_u64_1073_inst_req_0;
      CONCAT_u32_u64_1073_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u32_u64_1073_inst_req_1;
      CONCAT_u32_u64_1073_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_12_gI: SplitGuardInterface generic map(name => "ApConcat_group_12_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_12",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 12
    -- shared split operator group (13) : CONCAT_u32_u64_1099_inst 
    ApConcat_group_13: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u16_u32_1093_wire & CONCAT_u16_u32_1098_wire;
      CONCAT_u32_u64_1099_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u32_u64_1099_inst_req_0;
      CONCAT_u32_u64_1099_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u32_u64_1099_inst_req_1;
      CONCAT_u32_u64_1099_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_13_gI: SplitGuardInterface generic map(name => "ApConcat_group_13_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_13",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : CONCAT_u32_u64_1125_inst 
    ApConcat_group_14: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u16_u32_1119_wire & CONCAT_u16_u32_1124_wire;
      CONCAT_u32_u64_1125_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u32_u64_1125_inst_req_0;
      CONCAT_u32_u64_1125_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u32_u64_1125_inst_req_1;
      CONCAT_u32_u64_1125_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_14_gI: SplitGuardInterface generic map(name => "ApConcat_group_14_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_14",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- binary operator SGT_i16_u1_1004_inst
    process(a116_448, a216_512) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a116_448, a216_512, tmp_var);
      SGT_i16_u1_1004_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_1012_inst
    process(a316_576, a416_640) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a316_576, a416_640, tmp_var);
      SGT_i16_u1_1012_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_1020_inst
    process(t161_1008, t162_1016) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t161_1008, t162_1016, tmp_var);
      SGT_i16_u1_1020_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_644_inst
    process(a11_388, a21_452) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a11_388, a21_452, tmp_var);
      SGT_i16_u1_644_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_652_inst
    process(a31_516, a41_580) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a31_516, a41_580, tmp_var);
      SGT_i16_u1_652_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_660_inst
    process(t11_648, t12_656) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t11_648, t12_656, tmp_var);
      SGT_i16_u1_660_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_668_inst
    process(a12_392, a22_456) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a12_392, a22_456, tmp_var);
      SGT_i16_u1_668_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_676_inst
    process(a32_520, a42_584) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a32_520, a42_584, tmp_var);
      SGT_i16_u1_676_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_684_inst
    process(t21_672, t22_680) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t21_672, t22_680, tmp_var);
      SGT_i16_u1_684_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_692_inst
    process(a13_396, a23_460) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a13_396, a23_460, tmp_var);
      SGT_i16_u1_692_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_700_inst
    process(a33_524, a43_588) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a33_524, a43_588, tmp_var);
      SGT_i16_u1_700_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_708_inst
    process(t31_696, t32_704) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t31_696, t32_704, tmp_var);
      SGT_i16_u1_708_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_716_inst
    process(a14_400, a24_464) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a14_400, a24_464, tmp_var);
      SGT_i16_u1_716_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_724_inst
    process(a34_528, a44_592) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a34_528, a44_592, tmp_var);
      SGT_i16_u1_724_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_732_inst
    process(t41_720, t42_728) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t41_720, t42_728, tmp_var);
      SGT_i16_u1_732_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_740_inst
    process(a15_404, a25_468) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a15_404, a25_468, tmp_var);
      SGT_i16_u1_740_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_748_inst
    process(a35_532, a45_596) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a35_532, a45_596, tmp_var);
      SGT_i16_u1_748_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_756_inst
    process(t51_744, t52_752) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t51_744, t52_752, tmp_var);
      SGT_i16_u1_756_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_764_inst
    process(a16_408, a26_472) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a16_408, a26_472, tmp_var);
      SGT_i16_u1_764_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_772_inst
    process(a36_536, a46_600) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a36_536, a46_600, tmp_var);
      SGT_i16_u1_772_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_780_inst
    process(t61_768, t62_776) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t61_768, t62_776, tmp_var);
      SGT_i16_u1_780_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_788_inst
    process(a17_412, a27_476) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a17_412, a27_476, tmp_var);
      SGT_i16_u1_788_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_796_inst
    process(a37_540, a47_604) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a37_540, a47_604, tmp_var);
      SGT_i16_u1_796_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_804_inst
    process(t71_792, t72_800) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t71_792, t72_800, tmp_var);
      SGT_i16_u1_804_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_812_inst
    process(a18_416, a28_480) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a18_416, a28_480, tmp_var);
      SGT_i16_u1_812_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_820_inst
    process(a38_544, a48_608) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a38_544, a48_608, tmp_var);
      SGT_i16_u1_820_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_828_inst
    process(t81_816, t82_824) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t81_816, t82_824, tmp_var);
      SGT_i16_u1_828_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_836_inst
    process(a19_420, a29_484) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a19_420, a29_484, tmp_var);
      SGT_i16_u1_836_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_844_inst
    process(a39_548, a49_612) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a39_548, a49_612, tmp_var);
      SGT_i16_u1_844_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_852_inst
    process(t91_840, t92_848) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t91_840, t92_848, tmp_var);
      SGT_i16_u1_852_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_860_inst
    process(a110_424, a210_488) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a110_424, a210_488, tmp_var);
      SGT_i16_u1_860_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_868_inst
    process(a310_552, a410_616) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a310_552, a410_616, tmp_var);
      SGT_i16_u1_868_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_876_inst
    process(t101_864, t102_872) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t101_864, t102_872, tmp_var);
      SGT_i16_u1_876_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_884_inst
    process(a111_428, a211_492) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a111_428, a211_492, tmp_var);
      SGT_i16_u1_884_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_892_inst
    process(a311_556, a411_620) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a311_556, a411_620, tmp_var);
      SGT_i16_u1_892_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_900_inst
    process(t111_888, t112_896) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t111_888, t112_896, tmp_var);
      SGT_i16_u1_900_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_908_inst
    process(a112_432, a212_496) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a112_432, a212_496, tmp_var);
      SGT_i16_u1_908_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_916_inst
    process(a312_560, a412_624) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a312_560, a412_624, tmp_var);
      SGT_i16_u1_916_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_924_inst
    process(t121_912, t122_920) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t121_912, t122_920, tmp_var);
      SGT_i16_u1_924_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_932_inst
    process(a113_436, a213_500) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a113_436, a213_500, tmp_var);
      SGT_i16_u1_932_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_940_inst
    process(a313_564, a413_628) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a313_564, a413_628, tmp_var);
      SGT_i16_u1_940_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_948_inst
    process(t131_936, t132_944) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t131_936, t132_944, tmp_var);
      SGT_i16_u1_948_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_956_inst
    process(a114_440, a214_504) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a114_440, a214_504, tmp_var);
      SGT_i16_u1_956_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_964_inst
    process(a314_568, a414_632) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a314_568, a414_632, tmp_var);
      SGT_i16_u1_964_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_972_inst
    process(t141_960, t142_968) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t141_960, t142_968, tmp_var);
      SGT_i16_u1_972_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_980_inst
    process(a115_444, a215_508) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a115_444, a215_508, tmp_var);
      SGT_i16_u1_980_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_988_inst
    process(a315_572, a415_636) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a315_572, a415_636, tmp_var);
      SGT_i16_u1_988_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_996_inst
    process(t151_984, t152_992) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t151_984, t152_992, tmp_var);
      SGT_i16_u1_996_wire <= tmp_var; --
    end process;
    -- shared split operator group (63) : array_obj_ref_101_index_offset 
    ApIntAdd_group_63: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_addr3_100_scaled;
      array_obj_ref_101_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_101_index_offset_req_0;
      array_obj_ref_101_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_101_index_offset_req_1;
      array_obj_ref_101_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_63_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_63_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_63",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 63
    -- shared split operator group (64) : array_obj_ref_1029_index_offset 
    ApIntAdd_group_64: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_addr_1028_scaled;
      array_obj_ref_1029_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1029_index_offset_req_0;
      array_obj_ref_1029_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1029_index_offset_req_1;
      array_obj_ref_1029_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_64_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_64_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_64",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 64
    -- shared split operator group (65) : array_obj_ref_1055_index_offset 
    ApIntAdd_group_65: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ADD_u32_u32_1054_scaled;
      array_obj_ref_1055_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1055_index_offset_req_0;
      array_obj_ref_1055_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1055_index_offset_req_1;
      array_obj_ref_1055_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_65_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_65_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_65",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 65
    -- shared split operator group (66) : array_obj_ref_1081_index_offset 
    ApIntAdd_group_66: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ADD_u32_u32_1080_scaled;
      array_obj_ref_1081_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1081_index_offset_req_0;
      array_obj_ref_1081_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1081_index_offset_req_1;
      array_obj_ref_1081_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_66_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_66_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_66",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 66
    -- shared split operator group (67) : array_obj_ref_108_index_offset 
    ApIntAdd_group_67: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_addr4_107_scaled;
      array_obj_ref_108_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_108_index_offset_req_0;
      array_obj_ref_108_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_108_index_offset_req_1;
      array_obj_ref_108_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_67_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_67_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_67",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 67
    -- shared split operator group (68) : array_obj_ref_1107_index_offset 
    ApIntAdd_group_68: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ADD_u32_u32_1106_scaled;
      array_obj_ref_1107_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1107_index_offset_req_0;
      array_obj_ref_1107_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1107_index_offset_req_1;
      array_obj_ref_1107_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_68_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_68_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_68",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 68
    -- shared split operator group (69) : array_obj_ref_87_index_offset 
    ApIntAdd_group_69: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_addr1_86_scaled;
      array_obj_ref_87_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_87_index_offset_req_0;
      array_obj_ref_87_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_87_index_offset_req_1;
      array_obj_ref_87_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_69_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_69_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_69",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 69
    -- shared split operator group (70) : array_obj_ref_94_index_offset 
    ApIntAdd_group_70: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_addr2_93_scaled;
      array_obj_ref_94_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_94_index_offset_req_0;
      array_obj_ref_94_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_94_index_offset_req_1;
      array_obj_ref_94_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_70_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_70_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_70",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 70
    -- shared load operator group (0) : ptr_deref_113_load_0 ptr_deref_125_load_0 ptr_deref_117_load_0 ptr_deref_121_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(55 downto 0);
      signal data_out: std_logic_vector(1023 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 2, 2 => 2, 1 => 2, 0 => 2);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 2, 2 => 2, 1 => 2, 0 => 2);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 6, 1 => 6, 2 => 6, 3 => 6);
      -- 
    begin -- 
      reqL_unguarded(3) <= ptr_deref_113_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_125_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_117_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_121_load_0_req_0;
      ptr_deref_113_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_125_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_117_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_121_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= ptr_deref_113_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_125_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_117_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_121_load_0_req_1;
      ptr_deref_113_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_125_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_117_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_121_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_113_word_address_0 & ptr_deref_125_word_address_0 & ptr_deref_117_word_address_0 & ptr_deref_121_word_address_0;
      ptr_deref_113_data_0 <= data_out(1023 downto 768);
      ptr_deref_125_data_0 <= data_out(767 downto 512);
      ptr_deref_117_data_0 <= data_out(511 downto 256);
      ptr_deref_121_data_0 <= data_out(255 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 4,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 256,
        num_reqs => 4,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(255 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_1036_store_0 ptr_deref_1062_store_0 ptr_deref_1088_store_0 ptr_deref_1114_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(55 downto 0);
      signal data_in: std_logic_vector(255 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 2, 2 => 2, 1 => 2, 0 => 2);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 15, 2 => 15, 1 => 15, 0 => 15);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 6, 1 => 6, 2 => 6, 3 => 6);
      -- 
    begin -- 
      reqL_unguarded(3) <= ptr_deref_1036_store_0_req_0;
      reqL_unguarded(2) <= ptr_deref_1062_store_0_req_0;
      reqL_unguarded(1) <= ptr_deref_1088_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1114_store_0_req_0;
      ptr_deref_1036_store_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_1062_store_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_1088_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1114_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= ptr_deref_1036_store_0_req_1;
      reqR_unguarded(2) <= ptr_deref_1062_store_0_req_1;
      reqR_unguarded(1) <= ptr_deref_1088_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1114_store_0_req_1;
      ptr_deref_1036_store_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_1062_store_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_1088_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1114_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_3: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1036_word_address_0 & ptr_deref_1062_word_address_0 & ptr_deref_1088_word_address_0 & ptr_deref_1114_word_address_0;
      data_in <= ptr_deref_1036_data_0 & ptr_deref_1062_data_0 & ptr_deref_1088_data_0 & ptr_deref_1114_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 4,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 4,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end maxPool4_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity sendB is -- 
  generic (tag_length : integer); 
  port ( -- 
    size : in  std_logic_vector(31 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
    maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity sendB;
architecture sendB_arch of sendB is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal size_buffer :  std_logic_vector(31 downto 0);
  signal size_update_enable: Boolean;
  -- output port buffer signals
  signal sendB_CP_2125_start: Boolean;
  signal sendB_CP_2125_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_1248_inst_req_1 : boolean;
  signal addr_of_1198_final_reg_req_1 : boolean;
  signal if_stmt_1141_branch_ack_1 : boolean;
  signal type_cast_1248_inst_ack_1 : boolean;
  signal type_cast_1168_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1250_inst_req_0 : boolean;
  signal type_cast_1248_inst_req_0 : boolean;
  signal if_stmt_1141_branch_req_0 : boolean;
  signal type_cast_1248_inst_ack_0 : boolean;
  signal type_cast_1168_inst_req_1 : boolean;
  signal if_stmt_1141_branch_ack_0 : boolean;
  signal ptr_deref_1202_load_0_req_1 : boolean;
  signal addr_of_1198_final_reg_ack_1 : boolean;
  signal array_obj_ref_1197_index_offset_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1250_inst_ack_0 : boolean;
  signal array_obj_ref_1197_index_offset_req_1 : boolean;
  signal addr_of_1198_final_reg_ack_0 : boolean;
  signal ptr_deref_1202_load_0_ack_0 : boolean;
  signal array_obj_ref_1197_index_offset_ack_0 : boolean;
  signal array_obj_ref_1197_index_offset_req_0 : boolean;
  signal addr_of_1198_final_reg_req_0 : boolean;
  signal type_cast_1168_inst_req_0 : boolean;
  signal ptr_deref_1202_load_0_ack_1 : boolean;
  signal type_cast_1168_inst_ack_1 : boolean;
  signal type_cast_1255_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1257_inst_req_0 : boolean;
  signal type_cast_1255_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1257_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1257_inst_req_1 : boolean;
  signal type_cast_1255_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1250_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1250_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1257_inst_ack_1 : boolean;
  signal ptr_deref_1202_load_0_req_0 : boolean;
  signal type_cast_1255_inst_req_1 : boolean;
  signal type_cast_1262_inst_req_0 : boolean;
  signal type_cast_1262_inst_ack_0 : boolean;
  signal type_cast_1262_inst_req_1 : boolean;
  signal type_cast_1262_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1264_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1264_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1264_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1264_inst_ack_1 : boolean;
  signal type_cast_1269_inst_req_0 : boolean;
  signal type_cast_1269_inst_ack_0 : boolean;
  signal type_cast_1269_inst_req_1 : boolean;
  signal type_cast_1269_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1271_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1271_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1271_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1271_inst_ack_1 : boolean;
  signal type_cast_1276_inst_req_0 : boolean;
  signal type_cast_1276_inst_ack_0 : boolean;
  signal type_cast_1276_inst_req_1 : boolean;
  signal type_cast_1276_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1278_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1278_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1278_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1278_inst_ack_1 : boolean;
  signal type_cast_1283_inst_req_0 : boolean;
  signal type_cast_1283_inst_ack_0 : boolean;
  signal type_cast_1283_inst_req_1 : boolean;
  signal type_cast_1283_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1285_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1285_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1285_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1285_inst_ack_1 : boolean;
  signal type_cast_1290_inst_req_0 : boolean;
  signal type_cast_1290_inst_ack_0 : boolean;
  signal type_cast_1290_inst_req_1 : boolean;
  signal type_cast_1290_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1292_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1292_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1292_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1292_inst_ack_1 : boolean;
  signal type_cast_1297_inst_req_0 : boolean;
  signal type_cast_1297_inst_ack_0 : boolean;
  signal type_cast_1297_inst_req_1 : boolean;
  signal type_cast_1297_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1299_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1299_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1299_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1299_inst_ack_1 : boolean;
  signal if_stmt_1313_branch_req_0 : boolean;
  signal if_stmt_1313_branch_ack_1 : boolean;
  signal if_stmt_1313_branch_ack_0 : boolean;
  signal phi_stmt_1185_req_0 : boolean;
  signal type_cast_1191_inst_req_0 : boolean;
  signal type_cast_1191_inst_ack_0 : boolean;
  signal type_cast_1191_inst_req_1 : boolean;
  signal type_cast_1191_inst_ack_1 : boolean;
  signal phi_stmt_1185_req_1 : boolean;
  signal phi_stmt_1185_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "sendB_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 32) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= size;
  size_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(tag_length + 31 downto 32) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 31 downto 32);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  sendB_CP_2125_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "sendB_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendB_CP_2125_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sendB_CP_2125_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendB_CP_2125_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  sendB_CP_2125: Block -- control-path 
    signal sendB_CP_2125_elements: BooleanArray(59 downto 0);
    -- 
  begin -- 
    sendB_CP_2125_elements(0) <= sendB_CP_2125_start;
    sendB_CP_2125_symbol <= sendB_CP_2125_elements(59);
    -- CP-element group 0:  branch  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (15) 
      -- CP-element group 0: 	 branch_block_stmt_1134/assign_stmt_1140__entry__
      -- CP-element group 0: 	 branch_block_stmt_1134/assign_stmt_1140/$entry
      -- CP-element group 0: 	 branch_block_stmt_1134/if_stmt_1141_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_1134/assign_stmt_1140__exit__
      -- CP-element group 0: 	 branch_block_stmt_1134/R_cmp76_1142_place
      -- CP-element group 0: 	 branch_block_stmt_1134/if_stmt_1141__entry__
      -- CP-element group 0: 	 branch_block_stmt_1134/if_stmt_1141_if_link/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1134/assign_stmt_1140/$exit
      -- CP-element group 0: 	 branch_block_stmt_1134/if_stmt_1141_eval_test/branch_req
      -- CP-element group 0: 	 branch_block_stmt_1134/if_stmt_1141_eval_test/$entry
      -- CP-element group 0: 	 branch_block_stmt_1134/branch_block_stmt_1134__entry__
      -- CP-element group 0: 	 branch_block_stmt_1134/$entry
      -- CP-element group 0: 	 branch_block_stmt_1134/if_stmt_1141_else_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_1134/if_stmt_1141_eval_test/$exit
      -- 
    branch_req_2163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(0), ack => if_stmt_1141_branch_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	4 
    -- CP-element group 1: 	3 
    -- CP-element group 1:  members (18) 
      -- CP-element group 1: 	 branch_block_stmt_1134/if_stmt_1141_if_link/if_choice_transition
      -- CP-element group 1: 	 branch_block_stmt_1134/if_stmt_1141_if_link/$exit
      -- CP-element group 1: 	 branch_block_stmt_1134/assign_stmt_1153_to_assign_stmt_1182/type_cast_1168_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1134/entry_bbx_xnph
      -- CP-element group 1: 	 branch_block_stmt_1134/assign_stmt_1153_to_assign_stmt_1182/type_cast_1168_sample_start_
      -- CP-element group 1: 	 branch_block_stmt_1134/assign_stmt_1153_to_assign_stmt_1182/type_cast_1168_update_start_
      -- CP-element group 1: 	 branch_block_stmt_1134/merge_stmt_1147__exit__
      -- CP-element group 1: 	 branch_block_stmt_1134/assign_stmt_1153_to_assign_stmt_1182/type_cast_1168_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1134/assign_stmt_1153_to_assign_stmt_1182__entry__
      -- CP-element group 1: 	 branch_block_stmt_1134/assign_stmt_1153_to_assign_stmt_1182/type_cast_1168_Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1134/assign_stmt_1153_to_assign_stmt_1182/type_cast_1168_Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1134/assign_stmt_1153_to_assign_stmt_1182/$entry
      -- CP-element group 1: 	 branch_block_stmt_1134/entry_bbx_xnph_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_1134/entry_bbx_xnph_PhiReq/$exit
      -- CP-element group 1: 	 branch_block_stmt_1134/merge_stmt_1147_PhiReqMerge
      -- CP-element group 1: 	 branch_block_stmt_1134/merge_stmt_1147_PhiAck/$entry
      -- CP-element group 1: 	 branch_block_stmt_1134/merge_stmt_1147_PhiAck/$exit
      -- CP-element group 1: 	 branch_block_stmt_1134/merge_stmt_1147_PhiAck/dummy
      -- 
    if_choice_transition_2168_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1141_branch_ack_1, ack => sendB_CP_2125_elements(1)); -- 
    cr_2190_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2190_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(1), ack => type_cast_1168_inst_req_1); -- 
    rr_2185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(1), ack => type_cast_1168_inst_req_0); -- 
    -- CP-element group 2:  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	59 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 branch_block_stmt_1134/entry_forx_xend
      -- CP-element group 2: 	 branch_block_stmt_1134/if_stmt_1141_else_link/else_choice_transition
      -- CP-element group 2: 	 branch_block_stmt_1134/if_stmt_1141_else_link/$exit
      -- CP-element group 2: 	 branch_block_stmt_1134/entry_forx_xend_PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_1134/entry_forx_xend_PhiReq/$exit
      -- 
    else_choice_transition_2172_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1141_branch_ack_0, ack => sendB_CP_2125_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	1 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_1134/assign_stmt_1153_to_assign_stmt_1182/type_cast_1168_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1134/assign_stmt_1153_to_assign_stmt_1182/type_cast_1168_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_1134/assign_stmt_1153_to_assign_stmt_1182/type_cast_1168_Sample/$exit
      -- 
    ra_2186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1168_inst_ack_0, ack => sendB_CP_2125_elements(3)); -- 
    -- CP-element group 4:  transition  place  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	1 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	53 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_1134/assign_stmt_1153_to_assign_stmt_1182/$exit
      -- CP-element group 4: 	 branch_block_stmt_1134/assign_stmt_1153_to_assign_stmt_1182/type_cast_1168_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_1134/assign_stmt_1153_to_assign_stmt_1182__exit__
      -- CP-element group 4: 	 branch_block_stmt_1134/bbx_xnph_forx_xbody
      -- CP-element group 4: 	 branch_block_stmt_1134/assign_stmt_1153_to_assign_stmt_1182/type_cast_1168_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1134/assign_stmt_1153_to_assign_stmt_1182/type_cast_1168_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_1134/bbx_xnph_forx_xbody_PhiReq/$entry
      -- CP-element group 4: 	 branch_block_stmt_1134/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1185/$entry
      -- CP-element group 4: 	 branch_block_stmt_1134/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1185/phi_stmt_1185_sources/$entry
      -- 
    ca_2191_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1168_inst_ack_1, ack => sendB_CP_2125_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	58 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	50 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/array_obj_ref_1197_final_index_sum_regn_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/array_obj_ref_1197_final_index_sum_regn_sample_complete
      -- CP-element group 5: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/array_obj_ref_1197_final_index_sum_regn_Sample/ack
      -- 
    ack_2220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1197_index_offset_ack_0, ack => sendB_CP_2125_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	58 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (11) 
      -- CP-element group 6: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/addr_of_1198_request/$entry
      -- CP-element group 6: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/array_obj_ref_1197_offset_calculated
      -- CP-element group 6: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/array_obj_ref_1197_base_plus_offset/sum_rename_req
      -- CP-element group 6: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/array_obj_ref_1197_base_plus_offset/$exit
      -- CP-element group 6: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/array_obj_ref_1197_base_plus_offset/$entry
      -- CP-element group 6: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/array_obj_ref_1197_base_plus_offset/sum_rename_ack
      -- CP-element group 6: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/array_obj_ref_1197_final_index_sum_regn_Update/ack
      -- CP-element group 6: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/array_obj_ref_1197_final_index_sum_regn_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/array_obj_ref_1197_root_address_calculated
      -- CP-element group 6: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/addr_of_1198_request/req
      -- CP-element group 6: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/addr_of_1198_sample_start_
      -- 
    ack_2225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1197_index_offset_ack_1, ack => sendB_CP_2125_elements(6)); -- 
    req_2234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(6), ack => addr_of_1198_final_reg_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/addr_of_1198_request/$exit
      -- CP-element group 7: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/addr_of_1198_request/ack
      -- CP-element group 7: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/addr_of_1198_sample_completed_
      -- 
    ack_2235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1198_final_reg_ack_0, ack => sendB_CP_2125_elements(7)); -- 
    -- CP-element group 8:  join  fork  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	58 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (24) 
      -- CP-element group 8: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/ptr_deref_1202_base_address_resized
      -- CP-element group 8: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/ptr_deref_1202_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/addr_of_1198_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/addr_of_1198_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/ptr_deref_1202_word_addrgen/root_register_req
      -- CP-element group 8: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/ptr_deref_1202_word_addrgen/root_register_ack
      -- CP-element group 8: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/ptr_deref_1202_base_addr_resize/base_resize_ack
      -- CP-element group 8: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/ptr_deref_1202_base_addr_resize/$exit
      -- CP-element group 8: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/ptr_deref_1202_base_addr_resize/base_resize_req
      -- CP-element group 8: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/ptr_deref_1202_base_addr_resize/$entry
      -- CP-element group 8: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/ptr_deref_1202_base_plus_offset/$entry
      -- CP-element group 8: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/ptr_deref_1202_word_addrgen/$exit
      -- CP-element group 8: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/ptr_deref_1202_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/ptr_deref_1202_word_addrgen/$entry
      -- CP-element group 8: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/ptr_deref_1202_base_plus_offset/sum_rename_ack
      -- CP-element group 8: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/addr_of_1198_complete/ack
      -- CP-element group 8: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/ptr_deref_1202_base_plus_offset/sum_rename_req
      -- CP-element group 8: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/ptr_deref_1202_base_plus_offset/$exit
      -- CP-element group 8: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/ptr_deref_1202_Sample/word_access_start/$entry
      -- CP-element group 8: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/ptr_deref_1202_base_address_calculated
      -- CP-element group 8: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/ptr_deref_1202_Sample/word_access_start/word_0/$entry
      -- CP-element group 8: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/ptr_deref_1202_word_address_calculated
      -- CP-element group 8: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/ptr_deref_1202_Sample/word_access_start/word_0/rr
      -- CP-element group 8: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/ptr_deref_1202_root_address_calculated
      -- 
    ack_2240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1198_final_reg_ack_1, ack => sendB_CP_2125_elements(8)); -- 
    rr_2273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(8), ack => ptr_deref_1202_load_0_req_0); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/ptr_deref_1202_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/ptr_deref_1202_Sample/word_access_start/word_0/ra
      -- CP-element group 9: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/ptr_deref_1202_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/ptr_deref_1202_Sample/word_access_start/$exit
      -- CP-element group 9: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/ptr_deref_1202_Sample/word_access_start/word_0/$exit
      -- 
    ra_2274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1202_load_0_ack_0, ack => sendB_CP_2125_elements(9)); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	58 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	15 
    -- CP-element group 10: 	20 
    -- CP-element group 10: 	25 
    -- CP-element group 10: 	30 
    -- CP-element group 10: 	35 
    -- CP-element group 10: 	40 
    -- CP-element group 10: 	45 
    -- CP-element group 10:  members (33) 
      -- CP-element group 10: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/ptr_deref_1202_Update/word_access_complete/$exit
      -- CP-element group 10: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1248_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/ptr_deref_1202_Update/ptr_deref_1202_Merge/$entry
      -- CP-element group 10: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/ptr_deref_1202_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1248_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/ptr_deref_1202_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1248_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/ptr_deref_1202_Update/word_access_complete/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/ptr_deref_1202_Update/word_access_complete/word_0/ca
      -- CP-element group 10: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/ptr_deref_1202_Update/ptr_deref_1202_Merge/$exit
      -- CP-element group 10: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1255_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/ptr_deref_1202_Update/ptr_deref_1202_Merge/merge_req
      -- CP-element group 10: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1255_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1262_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1255_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/ptr_deref_1202_Update/ptr_deref_1202_Merge/merge_ack
      -- CP-element group 10: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1262_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1262_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1269_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1269_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1269_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1276_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1276_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1276_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1283_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1283_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1283_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1290_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1290_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1290_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1297_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1297_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1297_Sample/rr
      -- 
    ca_2285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1202_load_0_ack_1, ack => sendB_CP_2125_elements(10)); -- 
    rr_2298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(10), ack => type_cast_1248_inst_req_0); -- 
    rr_2326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(10), ack => type_cast_1255_inst_req_0); -- 
    rr_2354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(10), ack => type_cast_1262_inst_req_0); -- 
    rr_2382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(10), ack => type_cast_1269_inst_req_0); -- 
    rr_2410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(10), ack => type_cast_1276_inst_req_0); -- 
    rr_2438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(10), ack => type_cast_1283_inst_req_0); -- 
    rr_2466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(10), ack => type_cast_1290_inst_req_0); -- 
    rr_2494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(10), ack => type_cast_1297_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1248_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1248_Sample/ra
      -- CP-element group 11: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1248_sample_completed_
      -- 
    ra_2299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1248_inst_ack_0, ack => sendB_CP_2125_elements(11)); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	58 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1248_Update/ca
      -- CP-element group 12: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1248_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1250_Sample/req
      -- CP-element group 12: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1250_Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1250_sample_start_
      -- CP-element group 12: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1248_Update/$exit
      -- 
    ca_2304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1248_inst_ack_1, ack => sendB_CP_2125_elements(12)); -- 
    req_2312_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2312_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(12), ack => WPIPE_maxpool_output_pipe_1250_inst_req_0); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1250_Sample/ack
      -- CP-element group 13: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1250_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1250_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1250_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1250_Update/req
      -- CP-element group 13: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1250_update_start_
      -- 
    ack_2313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1250_inst_ack_0, ack => sendB_CP_2125_elements(13)); -- 
    req_2317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(13), ack => WPIPE_maxpool_output_pipe_1250_inst_req_1); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1250_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1250_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1250_Update/ack
      -- 
    ack_2318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1250_inst_ack_1, ack => sendB_CP_2125_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1255_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1255_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1255_sample_completed_
      -- 
    ra_2327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1255_inst_ack_0, ack => sendB_CP_2125_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	58 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1255_Update/ca
      -- CP-element group 16: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1255_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1255_Update/$exit
      -- 
    ca_2332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1255_inst_ack_1, ack => sendB_CP_2125_elements(16)); -- 
    -- CP-element group 17:  join  transition  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1257_Sample/req
      -- CP-element group 17: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1257_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1257_sample_start_
      -- 
    req_2340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(17), ack => WPIPE_maxpool_output_pipe_1257_inst_req_0); -- 
    sendB_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2125_elements(14) & sendB_CP_2125_elements(16);
      gj_sendB_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2125_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1257_Sample/ack
      -- CP-element group 18: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1257_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1257_Update/req
      -- CP-element group 18: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1257_update_start_
      -- CP-element group 18: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1257_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1257_sample_completed_
      -- 
    ack_2341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1257_inst_ack_0, ack => sendB_CP_2125_elements(18)); -- 
    req_2345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(18), ack => WPIPE_maxpool_output_pipe_1257_inst_req_1); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	22 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1257_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1257_Update/ack
      -- CP-element group 19: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1257_update_completed_
      -- 
    ack_2346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1257_inst_ack_1, ack => sendB_CP_2125_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	10 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1262_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1262_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1262_Sample/ra
      -- 
    ra_2355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1262_inst_ack_0, ack => sendB_CP_2125_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	58 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1262_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1262_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1262_Update/ca
      -- 
    ca_2360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1262_inst_ack_1, ack => sendB_CP_2125_elements(21)); -- 
    -- CP-element group 22:  join  transition  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	19 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1264_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1264_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1264_Sample/req
      -- 
    req_2368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(22), ack => WPIPE_maxpool_output_pipe_1264_inst_req_0); -- 
    sendB_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2125_elements(19) & sendB_CP_2125_elements(21);
      gj_sendB_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2125_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (6) 
      -- CP-element group 23: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1264_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1264_update_start_
      -- CP-element group 23: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1264_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1264_Sample/ack
      -- CP-element group 23: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1264_Update/$entry
      -- CP-element group 23: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1264_Update/req
      -- 
    ack_2369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1264_inst_ack_0, ack => sendB_CP_2125_elements(23)); -- 
    req_2373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(23), ack => WPIPE_maxpool_output_pipe_1264_inst_req_1); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	27 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1264_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1264_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1264_Update/ack
      -- 
    ack_2374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1264_inst_ack_1, ack => sendB_CP_2125_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	10 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1269_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1269_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1269_Sample/ra
      -- 
    ra_2383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1269_inst_ack_0, ack => sendB_CP_2125_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	58 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1269_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1269_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1269_Update/ca
      -- 
    ca_2388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1269_inst_ack_1, ack => sendB_CP_2125_elements(26)); -- 
    -- CP-element group 27:  join  transition  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	24 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1271_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1271_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1271_Sample/req
      -- 
    req_2396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(27), ack => WPIPE_maxpool_output_pipe_1271_inst_req_0); -- 
    sendB_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2125_elements(24) & sendB_CP_2125_elements(26);
      gj_sendB_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2125_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1271_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1271_update_start_
      -- CP-element group 28: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1271_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1271_Sample/ack
      -- CP-element group 28: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1271_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1271_Update/req
      -- 
    ack_2397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1271_inst_ack_0, ack => sendB_CP_2125_elements(28)); -- 
    req_2401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(28), ack => WPIPE_maxpool_output_pipe_1271_inst_req_1); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	32 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1271_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1271_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1271_Update/ack
      -- 
    ack_2402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1271_inst_ack_1, ack => sendB_CP_2125_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	10 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1276_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1276_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1276_Sample/ra
      -- 
    ra_2411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1276_inst_ack_0, ack => sendB_CP_2125_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	58 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1276_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1276_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1276_Update/ca
      -- 
    ca_2416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1276_inst_ack_1, ack => sendB_CP_2125_elements(31)); -- 
    -- CP-element group 32:  join  transition  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	29 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1278_sample_start_
      -- CP-element group 32: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1278_Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1278_Sample/req
      -- 
    req_2424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(32), ack => WPIPE_maxpool_output_pipe_1278_inst_req_0); -- 
    sendB_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2125_elements(29) & sendB_CP_2125_elements(31);
      gj_sendB_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2125_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1278_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1278_update_start_
      -- CP-element group 33: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1278_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1278_Sample/ack
      -- CP-element group 33: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1278_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1278_Update/req
      -- 
    ack_2425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1278_inst_ack_0, ack => sendB_CP_2125_elements(33)); -- 
    req_2429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(33), ack => WPIPE_maxpool_output_pipe_1278_inst_req_1); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	37 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1278_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1278_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1278_Update/ack
      -- 
    ack_2430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1278_inst_ack_1, ack => sendB_CP_2125_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	10 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1283_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1283_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1283_Sample/ra
      -- 
    ra_2439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1283_inst_ack_0, ack => sendB_CP_2125_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	58 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1283_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1283_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1283_Update/ca
      -- 
    ca_2444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1283_inst_ack_1, ack => sendB_CP_2125_elements(36)); -- 
    -- CP-element group 37:  join  transition  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1285_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1285_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1285_Sample/req
      -- 
    req_2452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(37), ack => WPIPE_maxpool_output_pipe_1285_inst_req_0); -- 
    sendB_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2125_elements(34) & sendB_CP_2125_elements(36);
      gj_sendB_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2125_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1285_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1285_update_start_
      -- CP-element group 38: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1285_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1285_Sample/ack
      -- CP-element group 38: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1285_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1285_Update/req
      -- 
    ack_2453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1285_inst_ack_0, ack => sendB_CP_2125_elements(38)); -- 
    req_2457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(38), ack => WPIPE_maxpool_output_pipe_1285_inst_req_1); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	42 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1285_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1285_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1285_Update/ack
      -- 
    ack_2458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1285_inst_ack_1, ack => sendB_CP_2125_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	10 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1290_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1290_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1290_Sample/ra
      -- 
    ra_2467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1290_inst_ack_0, ack => sendB_CP_2125_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	58 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1290_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1290_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1290_Update/ca
      -- 
    ca_2472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1290_inst_ack_1, ack => sendB_CP_2125_elements(41)); -- 
    -- CP-element group 42:  join  transition  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	39 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1292_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1292_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1292_Sample/req
      -- 
    req_2480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(42), ack => WPIPE_maxpool_output_pipe_1292_inst_req_0); -- 
    sendB_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2125_elements(39) & sendB_CP_2125_elements(41);
      gj_sendB_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2125_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (6) 
      -- CP-element group 43: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1292_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1292_update_start_
      -- CP-element group 43: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1292_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1292_Sample/ack
      -- CP-element group 43: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1292_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1292_Update/req
      -- 
    ack_2481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1292_inst_ack_0, ack => sendB_CP_2125_elements(43)); -- 
    req_2485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(43), ack => WPIPE_maxpool_output_pipe_1292_inst_req_1); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	47 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1292_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1292_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1292_Update/ack
      -- 
    ack_2486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1292_inst_ack_1, ack => sendB_CP_2125_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	10 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1297_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1297_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1297_Sample/ra
      -- 
    ra_2495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1297_inst_ack_0, ack => sendB_CP_2125_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	58 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1297_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1297_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1297_Update/ca
      -- 
    ca_2500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1297_inst_ack_1, ack => sendB_CP_2125_elements(46)); -- 
    -- CP-element group 47:  join  transition  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	44 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1299_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1299_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1299_Sample/req
      -- 
    req_2508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(47), ack => WPIPE_maxpool_output_pipe_1299_inst_req_0); -- 
    sendB_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2125_elements(44) & sendB_CP_2125_elements(46);
      gj_sendB_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2125_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (6) 
      -- CP-element group 48: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1299_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1299_update_start_
      -- CP-element group 48: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1299_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1299_Sample/ack
      -- CP-element group 48: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1299_Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1299_Update/req
      -- 
    ack_2509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1299_inst_ack_0, ack => sendB_CP_2125_elements(48)); -- 
    req_2513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(48), ack => WPIPE_maxpool_output_pipe_1299_inst_req_1); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1299_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1299_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/WPIPE_maxpool_output_pipe_1299_Update/ack
      -- 
    ack_2514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1299_inst_ack_1, ack => sendB_CP_2125_elements(49)); -- 
    -- CP-element group 50:  branch  join  transition  place  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	5 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (10) 
      -- CP-element group 50: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312__exit__
      -- CP-element group 50: 	 branch_block_stmt_1134/if_stmt_1313__entry__
      -- CP-element group 50: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/$exit
      -- CP-element group 50: 	 branch_block_stmt_1134/if_stmt_1313_dead_link/$entry
      -- CP-element group 50: 	 branch_block_stmt_1134/if_stmt_1313_eval_test/$entry
      -- CP-element group 50: 	 branch_block_stmt_1134/if_stmt_1313_eval_test/$exit
      -- CP-element group 50: 	 branch_block_stmt_1134/if_stmt_1313_eval_test/branch_req
      -- CP-element group 50: 	 branch_block_stmt_1134/R_exitcond1_1314_place
      -- CP-element group 50: 	 branch_block_stmt_1134/if_stmt_1313_if_link/$entry
      -- CP-element group 50: 	 branch_block_stmt_1134/if_stmt_1313_else_link/$entry
      -- 
    branch_req_2522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(50), ack => if_stmt_1313_branch_req_0); -- 
    sendB_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2125_elements(5) & sendB_CP_2125_elements(49);
      gj_sendB_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2125_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  merge  transition  place  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	59 
    -- CP-element group 51:  members (13) 
      -- CP-element group 51: 	 branch_block_stmt_1134/merge_stmt_1319__exit__
      -- CP-element group 51: 	 branch_block_stmt_1134/forx_xendx_xloopexit_forx_xend
      -- CP-element group 51: 	 branch_block_stmt_1134/if_stmt_1313_if_link/$exit
      -- CP-element group 51: 	 branch_block_stmt_1134/if_stmt_1313_if_link/if_choice_transition
      -- CP-element group 51: 	 branch_block_stmt_1134/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 51: 	 branch_block_stmt_1134/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 51: 	 branch_block_stmt_1134/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 51: 	 branch_block_stmt_1134/merge_stmt_1319_PhiReqMerge
      -- CP-element group 51: 	 branch_block_stmt_1134/merge_stmt_1319_PhiAck/$entry
      -- CP-element group 51: 	 branch_block_stmt_1134/merge_stmt_1319_PhiAck/$exit
      -- CP-element group 51: 	 branch_block_stmt_1134/merge_stmt_1319_PhiAck/dummy
      -- CP-element group 51: 	 branch_block_stmt_1134/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 51: 	 branch_block_stmt_1134/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_2527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1313_branch_ack_1, ack => sendB_CP_2125_elements(51)); -- 
    -- CP-element group 52:  fork  transition  place  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52: 	55 
    -- CP-element group 52:  members (12) 
      -- CP-element group 52: 	 branch_block_stmt_1134/if_stmt_1313_else_link/$exit
      -- CP-element group 52: 	 branch_block_stmt_1134/if_stmt_1313_else_link/else_choice_transition
      -- CP-element group 52: 	 branch_block_stmt_1134/forx_xbody_forx_xbody
      -- CP-element group 52: 	 branch_block_stmt_1134/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 52: 	 branch_block_stmt_1134/forx_xbody_forx_xbody_PhiReq/phi_stmt_1185/$entry
      -- CP-element group 52: 	 branch_block_stmt_1134/forx_xbody_forx_xbody_PhiReq/phi_stmt_1185/phi_stmt_1185_sources/$entry
      -- CP-element group 52: 	 branch_block_stmt_1134/forx_xbody_forx_xbody_PhiReq/phi_stmt_1185/phi_stmt_1185_sources/type_cast_1191/$entry
      -- CP-element group 52: 	 branch_block_stmt_1134/forx_xbody_forx_xbody_PhiReq/phi_stmt_1185/phi_stmt_1185_sources/type_cast_1191/SplitProtocol/$entry
      -- CP-element group 52: 	 branch_block_stmt_1134/forx_xbody_forx_xbody_PhiReq/phi_stmt_1185/phi_stmt_1185_sources/type_cast_1191/SplitProtocol/Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_1134/forx_xbody_forx_xbody_PhiReq/phi_stmt_1185/phi_stmt_1185_sources/type_cast_1191/SplitProtocol/Sample/rr
      -- CP-element group 52: 	 branch_block_stmt_1134/forx_xbody_forx_xbody_PhiReq/phi_stmt_1185/phi_stmt_1185_sources/type_cast_1191/SplitProtocol/Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_1134/forx_xbody_forx_xbody_PhiReq/phi_stmt_1185/phi_stmt_1185_sources/type_cast_1191/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1313_branch_ack_0, ack => sendB_CP_2125_elements(52)); -- 
    rr_2575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(52), ack => type_cast_1191_inst_req_0); -- 
    cr_2580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(52), ack => type_cast_1191_inst_req_1); -- 
    -- CP-element group 53:  transition  output  delay-element  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	4 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	57 
    -- CP-element group 53:  members (5) 
      -- CP-element group 53: 	 branch_block_stmt_1134/bbx_xnph_forx_xbody_PhiReq/$exit
      -- CP-element group 53: 	 branch_block_stmt_1134/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1185/$exit
      -- CP-element group 53: 	 branch_block_stmt_1134/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1185/phi_stmt_1185_sources/$exit
      -- CP-element group 53: 	 branch_block_stmt_1134/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1185/phi_stmt_1185_sources/type_cast_1189_konst_delay_trans
      -- CP-element group 53: 	 branch_block_stmt_1134/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1185/phi_stmt_1185_req
      -- 
    phi_stmt_1185_req_2556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1185_req_2556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(53), ack => phi_stmt_1185_req_0); -- 
    -- Element group sendB_CP_2125_elements(53) is a control-delay.
    cp_element_53_delay: control_delay_element  generic map(name => " 53_delay", delay_value => 1)  port map(req => sendB_CP_2125_elements(4), ack => sendB_CP_2125_elements(53), clk => clk, reset =>reset);
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (2) 
      -- CP-element group 54: 	 branch_block_stmt_1134/forx_xbody_forx_xbody_PhiReq/phi_stmt_1185/phi_stmt_1185_sources/type_cast_1191/SplitProtocol/Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_1134/forx_xbody_forx_xbody_PhiReq/phi_stmt_1185/phi_stmt_1185_sources/type_cast_1191/SplitProtocol/Sample/ra
      -- 
    ra_2576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1191_inst_ack_0, ack => sendB_CP_2125_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	52 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (2) 
      -- CP-element group 55: 	 branch_block_stmt_1134/forx_xbody_forx_xbody_PhiReq/phi_stmt_1185/phi_stmt_1185_sources/type_cast_1191/SplitProtocol/Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_1134/forx_xbody_forx_xbody_PhiReq/phi_stmt_1185/phi_stmt_1185_sources/type_cast_1191/SplitProtocol/Update/ca
      -- 
    ca_2581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1191_inst_ack_1, ack => sendB_CP_2125_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (6) 
      -- CP-element group 56: 	 branch_block_stmt_1134/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 56: 	 branch_block_stmt_1134/forx_xbody_forx_xbody_PhiReq/phi_stmt_1185/$exit
      -- CP-element group 56: 	 branch_block_stmt_1134/forx_xbody_forx_xbody_PhiReq/phi_stmt_1185/phi_stmt_1185_sources/$exit
      -- CP-element group 56: 	 branch_block_stmt_1134/forx_xbody_forx_xbody_PhiReq/phi_stmt_1185/phi_stmt_1185_sources/type_cast_1191/$exit
      -- CP-element group 56: 	 branch_block_stmt_1134/forx_xbody_forx_xbody_PhiReq/phi_stmt_1185/phi_stmt_1185_sources/type_cast_1191/SplitProtocol/$exit
      -- CP-element group 56: 	 branch_block_stmt_1134/forx_xbody_forx_xbody_PhiReq/phi_stmt_1185/phi_stmt_1185_req
      -- 
    phi_stmt_1185_req_2582_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1185_req_2582_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(56), ack => phi_stmt_1185_req_1); -- 
    sendB_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2125_elements(54) & sendB_CP_2125_elements(55);
      gj_sendB_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2125_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  merge  transition  place  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	53 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (2) 
      -- CP-element group 57: 	 branch_block_stmt_1134/merge_stmt_1184_PhiReqMerge
      -- CP-element group 57: 	 branch_block_stmt_1134/merge_stmt_1184_PhiAck/$entry
      -- 
    sendB_CP_2125_elements(57) <= OrReduce(sendB_CP_2125_elements(53) & sendB_CP_2125_elements(56));
    -- CP-element group 58:  fork  transition  place  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	12 
    -- CP-element group 58: 	16 
    -- CP-element group 58: 	5 
    -- CP-element group 58: 	6 
    -- CP-element group 58: 	8 
    -- CP-element group 58: 	10 
    -- CP-element group 58: 	21 
    -- CP-element group 58: 	26 
    -- CP-element group 58: 	31 
    -- CP-element group 58: 	36 
    -- CP-element group 58: 	41 
    -- CP-element group 58: 	46 
    -- CP-element group 58:  members (53) 
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1248_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/addr_of_1198_complete/req
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/ptr_deref_1202_Update/word_access_complete/word_0/$entry
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/array_obj_ref_1197_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/ptr_deref_1202_Update/word_access_complete/$entry
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/array_obj_ref_1197_final_index_sum_regn_update_start
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/array_obj_ref_1197_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/array_obj_ref_1197_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/ptr_deref_1202_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/ptr_deref_1202_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1248_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/array_obj_ref_1197_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/ptr_deref_1202_Update/word_access_complete/word_0/cr
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/array_obj_ref_1197_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/array_obj_ref_1197_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/array_obj_ref_1197_final_index_sum_regn_Update/req
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/array_obj_ref_1197_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/array_obj_ref_1197_final_index_sum_regn_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/array_obj_ref_1197_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/array_obj_ref_1197_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/array_obj_ref_1197_final_index_sum_regn_Sample/req
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/addr_of_1198_complete/$entry
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/array_obj_ref_1197_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/array_obj_ref_1197_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312__entry__
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1248_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/array_obj_ref_1197_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1134/merge_stmt_1184__exit__
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1262_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1255_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/$entry
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1255_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1255_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/addr_of_1198_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1262_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1262_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1269_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1269_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1269_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1276_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1276_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1276_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1283_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1283_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1283_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1290_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1290_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1290_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1297_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1297_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1134/assign_stmt_1199_to_assign_stmt_1312/type_cast_1297_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_1134/merge_stmt_1184_PhiAck/$exit
      -- CP-element group 58: 	 branch_block_stmt_1134/merge_stmt_1184_PhiAck/phi_stmt_1185_ack
      -- 
    phi_stmt_1185_ack_2587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1185_ack_0, ack => sendB_CP_2125_elements(58)); -- 
    cr_2303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(58), ack => type_cast_1248_inst_req_1); -- 
    req_2239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(58), ack => addr_of_1198_final_reg_req_1); -- 
    cr_2284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(58), ack => ptr_deref_1202_load_0_req_1); -- 
    req_2224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(58), ack => array_obj_ref_1197_index_offset_req_1); -- 
    req_2219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(58), ack => array_obj_ref_1197_index_offset_req_0); -- 
    cr_2331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(58), ack => type_cast_1255_inst_req_1); -- 
    cr_2359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(58), ack => type_cast_1262_inst_req_1); -- 
    cr_2387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(58), ack => type_cast_1269_inst_req_1); -- 
    cr_2415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(58), ack => type_cast_1276_inst_req_1); -- 
    cr_2443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(58), ack => type_cast_1283_inst_req_1); -- 
    cr_2471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(58), ack => type_cast_1290_inst_req_1); -- 
    cr_2499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2125_elements(58), ack => type_cast_1297_inst_req_1); -- 
    -- CP-element group 59:  merge  transition  place  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	2 
    -- CP-element group 59: 	51 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (16) 
      -- CP-element group 59: 	 branch_block_stmt_1134/merge_stmt_1323__exit__
      -- CP-element group 59: 	 $exit
      -- CP-element group 59: 	 branch_block_stmt_1134/$exit
      -- CP-element group 59: 	 branch_block_stmt_1134/branch_block_stmt_1134__exit__
      -- CP-element group 59: 	 branch_block_stmt_1134/merge_stmt_1321__exit__
      -- CP-element group 59: 	 branch_block_stmt_1134/return__
      -- CP-element group 59: 	 branch_block_stmt_1134/merge_stmt_1321_PhiReqMerge
      -- CP-element group 59: 	 branch_block_stmt_1134/merge_stmt_1321_PhiAck/$entry
      -- CP-element group 59: 	 branch_block_stmt_1134/merge_stmt_1321_PhiAck/$exit
      -- CP-element group 59: 	 branch_block_stmt_1134/merge_stmt_1321_PhiAck/dummy
      -- CP-element group 59: 	 branch_block_stmt_1134/return___PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_1134/return___PhiReq/$exit
      -- CP-element group 59: 	 branch_block_stmt_1134/merge_stmt_1323_PhiReqMerge
      -- CP-element group 59: 	 branch_block_stmt_1134/merge_stmt_1323_PhiAck/$entry
      -- CP-element group 59: 	 branch_block_stmt_1134/merge_stmt_1323_PhiAck/$exit
      -- CP-element group 59: 	 branch_block_stmt_1134/merge_stmt_1323_PhiAck/dummy
      -- 
    sendB_CP_2125_elements(59) <= OrReduce(sendB_CP_2125_elements(2) & sendB_CP_2125_elements(51));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar_1196_resized : std_logic_vector(13 downto 0);
    signal R_indvar_1196_scaled : std_logic_vector(13 downto 0);
    signal array_obj_ref_1197_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1197_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1197_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1197_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1197_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1197_root_address : std_logic_vector(13 downto 0);
    signal arrayidx_1199 : std_logic_vector(31 downto 0);
    signal cmp76_1140 : std_logic_vector(0 downto 0);
    signal conv52_1249 : std_logic_vector(7 downto 0);
    signal conv55_1256 : std_logic_vector(7 downto 0);
    signal conv58_1263 : std_logic_vector(7 downto 0);
    signal conv61_1270 : std_logic_vector(7 downto 0);
    signal conv64_1277 : std_logic_vector(7 downto 0);
    signal conv67_1284 : std_logic_vector(7 downto 0);
    signal conv70_1291 : std_logic_vector(7 downto 0);
    signal conv73_1298 : std_logic_vector(7 downto 0);
    signal exitcond1_1312 : std_logic_vector(0 downto 0);
    signal iNsTr_1_1169 : std_logic_vector(63 downto 0);
    signal indvar_1185 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1307 : std_logic_vector(63 downto 0);
    signal ptr_deref_1202_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1202_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1202_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1202_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1202_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr15_1215 : std_logic_vector(63 downto 0);
    signal shr21_1221 : std_logic_vector(63 downto 0);
    signal shr27_1227 : std_logic_vector(63 downto 0);
    signal shr33_1233 : std_logic_vector(63 downto 0);
    signal shr39_1239 : std_logic_vector(63 downto 0);
    signal shr45_1245 : std_logic_vector(63 downto 0);
    signal shr9_1209 : std_logic_vector(63 downto 0);
    signal shr_1153 : std_logic_vector(31 downto 0);
    signal shrx_xop_1165 : std_logic_vector(31 downto 0);
    signal tmp4_1203 : std_logic_vector(63 downto 0);
    signal tmp80_1182 : std_logic_vector(63 downto 0);
    signal tmp_1159 : std_logic_vector(0 downto 0);
    signal type_cast_1138_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1151_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1157_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1163_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1173_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1180_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1189_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1191_wire : std_logic_vector(63 downto 0);
    signal type_cast_1207_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1213_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1219_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1225_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1231_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1237_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1243_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1305_wire_constant : std_logic_vector(63 downto 0);
    signal xx_xop_1175 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1197_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1197_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1197_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1197_resized_base_address <= "00000000000000";
    ptr_deref_1202_word_offset_0 <= "00000000000000";
    type_cast_1138_wire_constant <= "00000000000000000000000000000011";
    type_cast_1151_wire_constant <= "00000000000000000000000000000010";
    type_cast_1157_wire_constant <= "00000000000000000000000000000001";
    type_cast_1163_wire_constant <= "11111111111111111111111111111111";
    type_cast_1173_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1180_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1189_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1207_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1213_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1219_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1225_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1231_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1237_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1243_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1305_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    phi_stmt_1185: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1189_wire_constant & type_cast_1191_wire;
      req <= phi_stmt_1185_req_0 & phi_stmt_1185_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1185",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1185_ack_0,
          idata => idata,
          odata => indvar_1185,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1185
    -- flow-through select operator MUX_1181_inst
    tmp80_1182 <= xx_xop_1175 when (tmp_1159(0) /=  '0') else type_cast_1180_wire_constant;
    addr_of_1198_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1198_final_reg_req_0;
      addr_of_1198_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1198_final_reg_req_1;
      addr_of_1198_final_reg_ack_1<= rack(0);
      addr_of_1198_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1198_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1197_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_1199,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1168_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1168_inst_req_0;
      type_cast_1168_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1168_inst_req_1;
      type_cast_1168_inst_ack_1<= rack(0);
      type_cast_1168_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1168_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shrx_xop_1165,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_1_1169,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1191_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1191_inst_req_0;
      type_cast_1191_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1191_inst_req_1;
      type_cast_1191_inst_ack_1<= rack(0);
      type_cast_1191_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1191_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1307,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1191_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1248_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1248_inst_req_0;
      type_cast_1248_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1248_inst_req_1;
      type_cast_1248_inst_ack_1<= rack(0);
      type_cast_1248_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1248_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr45_1245,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv52_1249,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1255_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1255_inst_req_0;
      type_cast_1255_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1255_inst_req_1;
      type_cast_1255_inst_ack_1<= rack(0);
      type_cast_1255_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1255_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr39_1239,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv55_1256,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1262_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1262_inst_req_0;
      type_cast_1262_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1262_inst_req_1;
      type_cast_1262_inst_ack_1<= rack(0);
      type_cast_1262_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1262_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr33_1233,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv58_1263,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1269_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1269_inst_req_0;
      type_cast_1269_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1269_inst_req_1;
      type_cast_1269_inst_ack_1<= rack(0);
      type_cast_1269_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1269_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr27_1227,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv61_1270,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1276_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1276_inst_req_0;
      type_cast_1276_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1276_inst_req_1;
      type_cast_1276_inst_ack_1<= rack(0);
      type_cast_1276_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1276_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr21_1221,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv64_1277,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1283_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1283_inst_req_0;
      type_cast_1283_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1283_inst_req_1;
      type_cast_1283_inst_ack_1<= rack(0);
      type_cast_1283_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1283_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr15_1215,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv67_1284,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1290_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1290_inst_req_0;
      type_cast_1290_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1290_inst_req_1;
      type_cast_1290_inst_ack_1<= rack(0);
      type_cast_1290_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1290_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr9_1209,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_1291,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1297_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1297_inst_req_0;
      type_cast_1297_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1297_inst_req_1;
      type_cast_1297_inst_ack_1<= rack(0);
      type_cast_1297_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1297_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp4_1203,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_1298,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1197_index_1_rename
    process(R_indvar_1196_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_1196_resized;
      ov(13 downto 0) := iv;
      R_indvar_1196_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1197_index_1_resize
    process(indvar_1185) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_1185;
      ov := iv(13 downto 0);
      R_indvar_1196_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1197_root_address_inst
    process(array_obj_ref_1197_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1197_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1197_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1202_addr_0
    process(ptr_deref_1202_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1202_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1202_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1202_base_resize
    process(arrayidx_1199) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_1199;
      ov := iv(13 downto 0);
      ptr_deref_1202_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1202_gather_scatter
    process(ptr_deref_1202_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1202_data_0;
      ov(63 downto 0) := iv;
      tmp4_1203 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1202_root_address_inst
    process(ptr_deref_1202_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1202_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1202_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1141_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp76_1140;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1141_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1141_branch_req_0,
          ack0 => if_stmt_1141_branch_ack_0,
          ack1 => if_stmt_1141_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1313_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_1312;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1313_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1313_branch_req_0,
          ack0 => if_stmt_1313_branch_ack_0,
          ack1 => if_stmt_1313_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_1164_inst
    process(shr_1153) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr_1153, type_cast_1163_wire_constant, tmp_var);
      shrx_xop_1165 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1174_inst
    process(iNsTr_1_1169) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_1_1169, type_cast_1173_wire_constant, tmp_var);
      xx_xop_1175 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1306_inst
    process(indvar_1185) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1185, type_cast_1305_wire_constant, tmp_var);
      indvarx_xnext_1307 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1311_inst
    process(indvarx_xnext_1307, tmp80_1182) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1307, tmp80_1182, tmp_var);
      exitcond1_1312 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1152_inst
    process(size_buffer) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(size_buffer, type_cast_1151_wire_constant, tmp_var);
      shr_1153 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1208_inst
    process(tmp4_1203) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_1203, type_cast_1207_wire_constant, tmp_var);
      shr9_1209 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1214_inst
    process(tmp4_1203) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_1203, type_cast_1213_wire_constant, tmp_var);
      shr15_1215 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1220_inst
    process(tmp4_1203) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_1203, type_cast_1219_wire_constant, tmp_var);
      shr21_1221 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1226_inst
    process(tmp4_1203) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_1203, type_cast_1225_wire_constant, tmp_var);
      shr27_1227 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1232_inst
    process(tmp4_1203) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_1203, type_cast_1231_wire_constant, tmp_var);
      shr33_1233 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1238_inst
    process(tmp4_1203) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_1203, type_cast_1237_wire_constant, tmp_var);
      shr39_1239 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1244_inst
    process(tmp4_1203) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_1203, type_cast_1243_wire_constant, tmp_var);
      shr45_1245 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1139_inst
    process(size_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(size_buffer, type_cast_1138_wire_constant, tmp_var);
      cmp76_1140 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1158_inst
    process(shr_1153) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(shr_1153, type_cast_1157_wire_constant, tmp_var);
      tmp_1159 <= tmp_var; --
    end process;
    -- shared split operator group (14) : array_obj_ref_1197_index_offset 
    ApIntAdd_group_14: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_1196_scaled;
      array_obj_ref_1197_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1197_index_offset_req_0;
      array_obj_ref_1197_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1197_index_offset_req_1;
      array_obj_ref_1197_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_14_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_14_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_14",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared load operator group (0) : ptr_deref_1202_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1202_load_0_req_0;
      ptr_deref_1202_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1202_load_0_req_1;
      ptr_deref_1202_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1202_word_address_0;
      ptr_deref_1202_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared outport operator group (0) : WPIPE_maxpool_output_pipe_1278_inst WPIPE_maxpool_output_pipe_1285_inst WPIPE_maxpool_output_pipe_1292_inst WPIPE_maxpool_output_pipe_1299_inst WPIPE_maxpool_output_pipe_1271_inst WPIPE_maxpool_output_pipe_1264_inst WPIPE_maxpool_output_pipe_1257_inst WPIPE_maxpool_output_pipe_1250_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 7 downto 0);
      signal update_req, update_ack : BooleanArray( 7 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 7 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      sample_req_unguarded(7) <= WPIPE_maxpool_output_pipe_1278_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_maxpool_output_pipe_1285_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_maxpool_output_pipe_1292_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_maxpool_output_pipe_1299_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_maxpool_output_pipe_1271_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_maxpool_output_pipe_1264_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1257_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1250_inst_req_0;
      WPIPE_maxpool_output_pipe_1278_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_maxpool_output_pipe_1285_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_maxpool_output_pipe_1292_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_maxpool_output_pipe_1299_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_maxpool_output_pipe_1271_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_1264_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_1257_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1250_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(7) <= WPIPE_maxpool_output_pipe_1278_inst_req_1;
      update_req_unguarded(6) <= WPIPE_maxpool_output_pipe_1285_inst_req_1;
      update_req_unguarded(5) <= WPIPE_maxpool_output_pipe_1292_inst_req_1;
      update_req_unguarded(4) <= WPIPE_maxpool_output_pipe_1299_inst_req_1;
      update_req_unguarded(3) <= WPIPE_maxpool_output_pipe_1271_inst_req_1;
      update_req_unguarded(2) <= WPIPE_maxpool_output_pipe_1264_inst_req_1;
      update_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1257_inst_req_1;
      update_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1250_inst_req_1;
      WPIPE_maxpool_output_pipe_1278_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_maxpool_output_pipe_1285_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_maxpool_output_pipe_1292_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_maxpool_output_pipe_1299_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_maxpool_output_pipe_1271_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_1264_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_1257_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1250_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      data_in <= conv64_1277 & conv67_1284 & conv70_1291 & conv73_1298 & conv61_1270 & conv58_1263 & conv55_1256 & conv52_1249;
      maxpool_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "maxpool_output_pipe_write_0_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      maxpool_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "maxpool_output_pipe", data_width => 8, num_reqs => 8, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => maxpool_output_pipe_pipe_write_req(0),
          oack => maxpool_output_pipe_pipe_write_ack(0),
          odata => maxpool_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end sendB_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    maxpool_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    maxpool_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    maxpool_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(19 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(2 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(2 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(19 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(255 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(2 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(255 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(2 downto 0);
  -- declarations related to module fill_T
  component fill_T is -- 
    generic (tag_length : integer); 
    port ( -- 
      addr : in  std_logic_vector(63 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(255 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(2 downto 0);
      maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module fill_T
  signal fill_T_addr :  std_logic_vector(63 downto 0);
  signal fill_T_in_args    : std_logic_vector(63 downto 0);
  signal fill_T_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal fill_T_tag_out   : std_logic_vector(1 downto 0);
  signal fill_T_start_req : std_logic;
  signal fill_T_start_ack : std_logic;
  signal fill_T_fin_req   : std_logic;
  signal fill_T_fin_ack : std_logic;
  -- caller side aggregated signals for module fill_T
  signal fill_T_call_reqs: std_logic_vector(0 downto 0);
  signal fill_T_call_acks: std_logic_vector(0 downto 0);
  signal fill_T_return_reqs: std_logic_vector(0 downto 0);
  signal fill_T_return_acks: std_logic_vector(0 downto 0);
  signal fill_T_call_data: std_logic_vector(63 downto 0);
  signal fill_T_call_tag: std_logic_vector(0 downto 0);
  signal fill_T_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module maxPool3D
  component maxPool3D is -- 
    generic (tag_length : integer); 
    port ( -- 
      maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      fill_T_call_reqs : out  std_logic_vector(0 downto 0);
      fill_T_call_acks : in   std_logic_vector(0 downto 0);
      fill_T_call_data : out  std_logic_vector(63 downto 0);
      fill_T_call_tag  :  out  std_logic_vector(0 downto 0);
      fill_T_return_reqs : out  std_logic_vector(0 downto 0);
      fill_T_return_acks : in   std_logic_vector(0 downto 0);
      fill_T_return_tag :  in   std_logic_vector(0 downto 0);
      maxPool4_call_reqs : out  std_logic_vector(0 downto 0);
      maxPool4_call_acks : in   std_logic_vector(0 downto 0);
      maxPool4_call_data : out  std_logic_vector(159 downto 0);
      maxPool4_call_tag  :  out  std_logic_vector(0 downto 0);
      maxPool4_return_reqs : out  std_logic_vector(0 downto 0);
      maxPool4_return_acks : in   std_logic_vector(0 downto 0);
      maxPool4_return_data : in   std_logic_vector(7 downto 0);
      maxPool4_return_tag :  in   std_logic_vector(0 downto 0);
      sendB_call_reqs : out  std_logic_vector(0 downto 0);
      sendB_call_acks : in   std_logic_vector(0 downto 0);
      sendB_call_data : out  std_logic_vector(31 downto 0);
      sendB_call_tag  :  out  std_logic_vector(0 downto 0);
      sendB_return_reqs : out  std_logic_vector(0 downto 0);
      sendB_return_acks : in   std_logic_vector(0 downto 0);
      sendB_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module maxPool3D
  signal maxPool3D_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal maxPool3D_tag_out   : std_logic_vector(1 downto 0);
  signal maxPool3D_start_req : std_logic;
  signal maxPool3D_start_ack : std_logic;
  signal maxPool3D_fin_req   : std_logic;
  signal maxPool3D_fin_ack : std_logic;
  -- declarations related to module maxPool4
  component maxPool4 is -- 
    generic (tag_length : integer); 
    port ( -- 
      addr : in  std_logic_vector(31 downto 0);
      addr1 : in  std_logic_vector(31 downto 0);
      addr2 : in  std_logic_vector(31 downto 0);
      addr3 : in  std_logic_vector(31 downto 0);
      addr4 : in  std_logic_vector(31 downto 0);
      output : out  std_logic_vector(7 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(255 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module maxPool4
  signal maxPool4_addr :  std_logic_vector(31 downto 0);
  signal maxPool4_addr1 :  std_logic_vector(31 downto 0);
  signal maxPool4_addr2 :  std_logic_vector(31 downto 0);
  signal maxPool4_addr3 :  std_logic_vector(31 downto 0);
  signal maxPool4_addr4 :  std_logic_vector(31 downto 0);
  signal maxPool4_output :  std_logic_vector(7 downto 0);
  signal maxPool4_in_args    : std_logic_vector(159 downto 0);
  signal maxPool4_out_args   : std_logic_vector(7 downto 0);
  signal maxPool4_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal maxPool4_tag_out   : std_logic_vector(1 downto 0);
  signal maxPool4_start_req : std_logic;
  signal maxPool4_start_ack : std_logic;
  signal maxPool4_fin_req   : std_logic;
  signal maxPool4_fin_ack : std_logic;
  -- caller side aggregated signals for module maxPool4
  signal maxPool4_call_reqs: std_logic_vector(0 downto 0);
  signal maxPool4_call_acks: std_logic_vector(0 downto 0);
  signal maxPool4_return_reqs: std_logic_vector(0 downto 0);
  signal maxPool4_return_acks: std_logic_vector(0 downto 0);
  signal maxPool4_call_data: std_logic_vector(159 downto 0);
  signal maxPool4_call_tag: std_logic_vector(0 downto 0);
  signal maxPool4_return_data: std_logic_vector(7 downto 0);
  signal maxPool4_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module sendB
  component sendB is -- 
    generic (tag_length : integer); 
    port ( -- 
      size : in  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module sendB
  signal sendB_size :  std_logic_vector(31 downto 0);
  signal sendB_in_args    : std_logic_vector(31 downto 0);
  signal sendB_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal sendB_tag_out   : std_logic_vector(1 downto 0);
  signal sendB_start_req : std_logic;
  signal sendB_start_ack : std_logic;
  signal sendB_fin_req   : std_logic;
  signal sendB_fin_ack : std_logic;
  -- caller side aggregated signals for module sendB
  signal sendB_call_reqs: std_logic_vector(0 downto 0);
  signal sendB_call_acks: std_logic_vector(0 downto 0);
  signal sendB_return_reqs: std_logic_vector(0 downto 0);
  signal sendB_return_acks: std_logic_vector(0 downto 0);
  signal sendB_call_data: std_logic_vector(31 downto 0);
  signal sendB_call_tag: std_logic_vector(0 downto 0);
  signal sendB_return_tag: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe maxpool_input_pipe
  signal maxpool_input_pipe_pipe_read_data: std_logic_vector(15 downto 0);
  signal maxpool_input_pipe_pipe_read_req: std_logic_vector(1 downto 0);
  signal maxpool_input_pipe_pipe_read_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe maxpool_output_pipe
  signal maxpool_output_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal maxpool_output_pipe_pipe_write_req: std_logic_vector(1 downto 0);
  signal maxpool_output_pipe_pipe_write_ack: std_logic_vector(1 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module fill_T
  fill_T_addr <= fill_T_in_args(63 downto 0);
  -- call arbiter for module fill_T
  fill_T_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => fill_T_call_reqs,
      call_acks => fill_T_call_acks,
      return_reqs => fill_T_return_reqs,
      return_acks => fill_T_return_acks,
      call_data  => fill_T_call_data,
      call_tag  => fill_T_call_tag,
      return_tag  => fill_T_return_tag,
      call_mtag => fill_T_tag_in,
      return_mtag => fill_T_tag_out,
      call_mreq => fill_T_start_req,
      call_mack => fill_T_start_ack,
      return_mreq => fill_T_fin_req,
      return_mack => fill_T_fin_ack,
      call_mdata => fill_T_in_args,
      clk => clk, 
      reset => reset --
    ); --
  fill_T_instance:fill_T-- 
    generic map(tag_length => 2)
    port map(-- 
      addr => fill_T_addr,
      start_req => fill_T_start_req,
      start_ack => fill_T_start_ack,
      fin_req => fill_T_fin_req,
      fin_ack => fill_T_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(255 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(19 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(2 downto 0),
      maxpool_input_pipe_pipe_read_req => maxpool_input_pipe_pipe_read_req(1 downto 1),
      maxpool_input_pipe_pipe_read_ack => maxpool_input_pipe_pipe_read_ack(1 downto 1),
      maxpool_input_pipe_pipe_read_data => maxpool_input_pipe_pipe_read_data(15 downto 8),
      tag_in => fill_T_tag_in,
      tag_out => fill_T_tag_out-- 
    ); -- 
  -- module maxPool3D
  maxPool3D_instance:maxPool3D-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => maxPool3D_start_req,
      start_ack => maxPool3D_start_ack,
      fin_req => maxPool3D_fin_req,
      fin_ack => maxPool3D_fin_ack,
      clk => clk,
      reset => reset,
      maxpool_input_pipe_pipe_read_req => maxpool_input_pipe_pipe_read_req(0 downto 0),
      maxpool_input_pipe_pipe_read_ack => maxpool_input_pipe_pipe_read_ack(0 downto 0),
      maxpool_input_pipe_pipe_read_data => maxpool_input_pipe_pipe_read_data(7 downto 0),
      maxpool_output_pipe_pipe_write_req => maxpool_output_pipe_pipe_write_req(0 downto 0),
      maxpool_output_pipe_pipe_write_ack => maxpool_output_pipe_pipe_write_ack(0 downto 0),
      maxpool_output_pipe_pipe_write_data => maxpool_output_pipe_pipe_write_data(7 downto 0),
      fill_T_call_reqs => fill_T_call_reqs(0 downto 0),
      fill_T_call_acks => fill_T_call_acks(0 downto 0),
      fill_T_call_data => fill_T_call_data(63 downto 0),
      fill_T_call_tag => fill_T_call_tag(0 downto 0),
      fill_T_return_reqs => fill_T_return_reqs(0 downto 0),
      fill_T_return_acks => fill_T_return_acks(0 downto 0),
      fill_T_return_tag => fill_T_return_tag(0 downto 0),
      maxPool4_call_reqs => maxPool4_call_reqs(0 downto 0),
      maxPool4_call_acks => maxPool4_call_acks(0 downto 0),
      maxPool4_call_data => maxPool4_call_data(159 downto 0),
      maxPool4_call_tag => maxPool4_call_tag(0 downto 0),
      maxPool4_return_reqs => maxPool4_return_reqs(0 downto 0),
      maxPool4_return_acks => maxPool4_return_acks(0 downto 0),
      maxPool4_return_data => maxPool4_return_data(7 downto 0),
      maxPool4_return_tag => maxPool4_return_tag(0 downto 0),
      sendB_call_reqs => sendB_call_reqs(0 downto 0),
      sendB_call_acks => sendB_call_acks(0 downto 0),
      sendB_call_data => sendB_call_data(31 downto 0),
      sendB_call_tag => sendB_call_tag(0 downto 0),
      sendB_return_reqs => sendB_return_reqs(0 downto 0),
      sendB_return_acks => sendB_return_acks(0 downto 0),
      sendB_return_tag => sendB_return_tag(0 downto 0),
      tag_in => maxPool3D_tag_in,
      tag_out => maxPool3D_tag_out-- 
    ); -- 
  -- module will be run forever 
  maxPool3D_tag_in <= (others => '0');
  maxPool3D_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => maxPool3D_start_req, start_ack => maxPool3D_start_ack,  fin_req => maxPool3D_fin_req,  fin_ack => maxPool3D_fin_ack);
  -- module maxPool4
  maxPool4_addr <= maxPool4_in_args(159 downto 128);
  maxPool4_addr1 <= maxPool4_in_args(127 downto 96);
  maxPool4_addr2 <= maxPool4_in_args(95 downto 64);
  maxPool4_addr3 <= maxPool4_in_args(63 downto 32);
  maxPool4_addr4 <= maxPool4_in_args(31 downto 0);
  maxPool4_out_args <= maxPool4_output ;
  -- call arbiter for module maxPool4
  maxPool4_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 160,
      return_data_width => 8,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => maxPool4_call_reqs,
      call_acks => maxPool4_call_acks,
      return_reqs => maxPool4_return_reqs,
      return_acks => maxPool4_return_acks,
      call_data  => maxPool4_call_data,
      call_tag  => maxPool4_call_tag,
      return_tag  => maxPool4_return_tag,
      call_mtag => maxPool4_tag_in,
      return_mtag => maxPool4_tag_out,
      return_data =>maxPool4_return_data,
      call_mreq => maxPool4_start_req,
      call_mack => maxPool4_start_ack,
      return_mreq => maxPool4_fin_req,
      return_mack => maxPool4_fin_ack,
      call_mdata => maxPool4_in_args,
      return_mdata => maxPool4_out_args,
      clk => clk, 
      reset => reset --
    ); --
  maxPool4_instance:maxPool4-- 
    generic map(tag_length => 2)
    port map(-- 
      addr => maxPool4_addr,
      addr1 => maxPool4_addr1,
      addr2 => maxPool4_addr2,
      addr3 => maxPool4_addr3,
      addr4 => maxPool4_addr4,
      output => maxPool4_output,
      start_req => maxPool4_start_req,
      start_ack => maxPool4_start_ack,
      fin_req => maxPool4_fin_req,
      fin_ack => maxPool4_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(19 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(255 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(2 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(13 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(19 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(2 downto 0),
      tag_in => maxPool4_tag_in,
      tag_out => maxPool4_tag_out-- 
    ); -- 
  -- module sendB
  sendB_size <= sendB_in_args(31 downto 0);
  -- call arbiter for module sendB
  sendB_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 32,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => sendB_call_reqs,
      call_acks => sendB_call_acks,
      return_reqs => sendB_return_reqs,
      return_acks => sendB_return_acks,
      call_data  => sendB_call_data,
      call_tag  => sendB_call_tag,
      return_tag  => sendB_return_tag,
      call_mtag => sendB_tag_in,
      return_mtag => sendB_tag_out,
      call_mreq => sendB_start_req,
      call_mack => sendB_start_ack,
      return_mreq => sendB_fin_req,
      return_mack => sendB_fin_ack,
      call_mdata => sendB_in_args,
      clk => clk, 
      reset => reset --
    ); --
  sendB_instance:sendB-- 
    generic map(tag_length => 2)
    port map(-- 
      size => sendB_size,
      start_req => sendB_start_req,
      start_ack => sendB_start_ack,
      fin_req => sendB_fin_req,
      fin_ack => sendB_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(19 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(2 downto 0),
      maxpool_output_pipe_pipe_write_req => maxpool_output_pipe_pipe_write_req(1 downto 1),
      maxpool_output_pipe_pipe_write_ack => maxpool_output_pipe_pipe_write_ack(1 downto 1),
      maxpool_output_pipe_pipe_write_data => maxpool_output_pipe_pipe_write_data(15 downto 8),
      tag_in => sendB_tag_in,
      tag_out => sendB_tag_out-- 
    ); -- 
  maxpool_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe maxpool_input_pipe",
      num_reads => 2,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => maxpool_input_pipe_pipe_read_req,
      read_ack => maxpool_input_pipe_pipe_read_ack,
      read_data => maxpool_input_pipe_pipe_read_data,
      write_req => maxpool_input_pipe_pipe_write_req,
      write_ack => maxpool_input_pipe_pipe_write_ack,
      write_data => maxpool_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  maxpool_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe maxpool_output_pipe",
      num_reads => 1,
      num_writes => 2,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => maxpool_output_pipe_pipe_read_req,
      read_ack => maxpool_output_pipe_pipe_read_ack,
      read_data => maxpool_output_pipe_pipe_read_data,
      write_req => maxpool_output_pipe_pipe_write_req,
      write_ack => maxpool_output_pipe_pipe_write_ack,
      write_data => maxpool_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 3,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 256,
      tag_width => 3,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 256
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
